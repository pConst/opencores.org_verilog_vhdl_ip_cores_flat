000000 => x"bc05", -- B
000001 => x"bc00", -- B
000002 => x"bc00", -- B
000003 => x"bc00", -- B
000004 => x"bc00", -- B
000005 => x"2800", -- CLR
000006 => x"ed0f", -- MCR
000007 => x"c2b2", -- LDIL
000008 => x"be09", -- BL
000009 => x"ed0f", -- MCR
000010 => x"3c00", -- SFT
000011 => x"0001", -- INC
000012 => x"c08f", -- LDIL
000013 => x"2001", -- AND
000014 => x"3c00", -- SFT
000015 => x"ed0f", -- MCR
000016 => x"bdf7", -- B
000017 => x"c77f", -- LDIL
000018 => x"0769", -- DECS
000019 => x"85ff", -- BNE
000020 => x"06d9", -- DECS
000021 => x"85fc", -- BNE
000022 => x"3470", -- RET
others => x"0000"  -- NOP