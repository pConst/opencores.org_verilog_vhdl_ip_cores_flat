// *****************************************************************************************
// 
// Version 0.2
// Modified 17.06.2007
// Designed by Ruslan Lepetenok
// *****************************************************************************************

// package tech_def_pack is

localparam c_tech_generic     = 0;

// Xilinx
localparam c_tech_virtex      = 1;
localparam c_tech_virtex_e    = 2;
localparam c_tech_virtex_ii   = 3;
localparam c_tech_virtex_4    = 4;
localparam c_tech_virtex_5    = 5; 
localparam c_tech_spartan_3   = 6;

// Altera
localparam c_tech_acex             = 7;

// end tech_def_pack;	
	
	
