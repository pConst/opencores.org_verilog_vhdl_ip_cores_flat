-------------------------------------------------------------------------------
-- Title: Serially Programmable Clock Source ICS307
-- Project: FH-Hagenberg/HSSE: SET5
-- Author: Copyright 2006 by Friedrich Seebacher and Markus Pfaff,
-- Linz/Austria/Europe
-------------------------------------------------------------------------------
-- $LastChangedDate: 2007-01-09 08:40:02 +0100 (Di, 09 Jän 2007) $
-- $LastChangedRevision: 415 $
-- $LastChangedBy: pfaff $
-- $HeadURL: file:///C:/pfaff/rpySvn/rpySvnSet5/trunk/Uebung/W06Jg04/Uebung03/unitIcs307/src/ICS307-e.vhd $
-- LoginNames: pfaff - Markus Pfaff, Linz/Austria/Europe
-------------------------------------------------------------------------------
-- Description: This description mimics a subset of the behaviour of the ICS307-02
-- versatile serially programmable clock source. This device is used as main clock
-- source on the SandboxX rapid prototyping system in HSSE and ESD courses at
-- FH-OOe/Hagenberg.
-- Due to the limited resolution of VHDL simulators when not used with fs as smallest
-- grain of time the unit will not transition frequency in the smooth way you'll read from
-- the data sheet. Instead it will transition from the old frequency value to the new one
-- after the transitioning time is over in a few steps.
-- Transitioning will get smoother with smaller transition times (gClkFrequcenyTransitionTime).
-- A transition time of several microseconds is not realistic, but will lead to a smooth
-- transition in simulation even if the simulator is set to ps resolution.
-- If time resolution is set to the minimum value (1 fs) you'll see a nice 
-- linear transition from one frequency to the other in your simulation.
-------------------------------------------------------------------------------
-- Not tested:
-- - Reconfiguring the ICS to a new frequency while the device is still transitioning.
-- - Reconfiguring the ICS several times
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ICS307 is
  generic (
    gInputFrequency             : natural := 25E6;  -- Reference input clock frequency [Hz]
    gClkFrequcenyTransitionTime : time    := 3 ms);

  port (
    -- SPI clock input
    iSclk   : in  std_ulogic;
    -- SPI data input
    iData   : in  std_ulogic;
    -- SPI strobe: latch data on falling edge of this signal
    iStrobe : in  std_ulogic;
    -- Clock signal generated by this unit
    oClk1   : out std_ulogic
    );
end ICS307;
