-- obj_code_pkg -- Object code in VHDL constant table for BRAM initialization.
-- Generated automatically with script 'build_rom.py'.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.l80pkg.all;

package obj_code_pkg is

constant obj_code : obj_code_t(0 to 313) := (
    X"c3", X"60", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c6", X"01", X"fb", X"c9", X"00", X"00", X"00", X"00", 
    X"3c", X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"3c", X"00", X"00", X"00", X"ef", X"00", X"00", X"00", 
    X"23", X"00", X"00", X"00", X"3e", X"42", X"00", X"00", 
    X"21", X"34", X"12", X"00", X"c3", X"2f", X"01", X"00", 
    X"cd", X"34", X"01", X"00", X"cd", X"37", X"01", X"00", 
    X"31", X"7a", X"01", X"3e", X"13", X"e7", X"fe", X"14", 
    X"c2", X"2a", X"01", X"3e", X"00", X"d3", X"10", X"fb", 
    X"3e", X"14", X"d3", X"11", X"3e", X"27", X"00", X"00", 
    X"00", X"00", X"fe", X"28", X"c2", X"2a", X"01", X"3e", 
    X"01", X"d3", X"10", X"fb", X"3e", X"14", X"d3", X"11", 
    X"3e", X"20", X"00", X"00", X"00", X"00", X"fe", X"21", 
    X"c2", X"2a", X"01", X"21", X"ff", X"13", X"3e", X"02", 
    X"d3", X"10", X"fb", X"3e", X"04", X"d3", X"11", X"00", 
    X"00", X"7d", X"fe", X"00", X"c2", X"2a", X"01", X"7c", 
    X"fe", X"14", X"c2", X"2a", X"01", X"3e", X"03", X"d3", 
    X"10", X"fb", X"3e", X"04", X"d3", X"11", X"00", X"00", 
    X"fe", X"42", X"c2", X"2a", X"01", X"3e", X"04", X"d3", 
    X"10", X"fb", X"3e", X"04", X"d3", X"11", X"00", X"00", 
    X"7c", X"fe", X"12", X"c2", X"2a", X"01", X"7d", X"fe", 
    X"34", X"c2", X"2a", X"01", X"3e", X"05", X"d3", X"10", 
    X"fb", X"3e", X"04", X"d3", X"11", X"00", X"00", X"fe", 
    X"79", X"c2", X"2a", X"01", X"3e", X"06", X"d3", X"10", 
    X"fb", X"3e", X"04", X"d3", X"11", X"3c", X"00", X"fe", 
    X"05", X"c2", X"2a", X"01", X"78", X"fe", X"19", X"c2", 
    X"2a", X"01", X"f3", X"3e", X"07", X"d3", X"10", X"3e", 
    X"04", X"d3", X"11", X"00", X"00", X"00", X"3e", X"50", 
    X"d3", X"12", X"3e", X"01", X"d3", X"10", X"fb", X"3e", 
    X"14", X"d3", X"11", X"3e", X"27", X"00", X"00", X"3c", 
    X"00", X"00", X"3c", X"00", X"00", X"00", X"00", X"00", 
    X"fe", X"2b", X"c2", X"2a", X"01", X"3e", X"55", X"d3", 
    X"20", X"76", X"3e", X"aa", X"d3", X"20", X"76", X"3e", 
    X"79", X"c3", X"df", X"00", X"06", X"19", X"c9", X"c3", 
    X"2a", X"01" 
);

end package obj_code_pkg;
