-- This is a block of initialized BRAM that contains the whole 4K Altair basic
-- image upon startup. The program starts at address zero so upon reset the
-- CPU will enter the 4K Basic code exactly as if it had been loaded from 
-- external media.
-- If the code in this block ever becomes corrupt, the only way to restore it
-- is reloading the FPGA.
-- This memory block is RAM; actually, it all the RAM the 4K demo needs to run.
-- The ROM identifiers below are a leftover from a previous version.


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity c2sb_4kbasic_rom is
    port ( 
        clk           : in std_logic;
        addr          : in std_logic_vector(15 downto 0);
        we            : in std_logic;
        data_in       : in std_logic_vector(7 downto 0);
        data_out      : out std_logic_vector(7 downto 0)
    );
end c2sb_4kbasic_rom;

architecture internal of c2sb_4kbasic_rom is

signal rom_addr :         std_logic_vector(11 downto 0);
type t_rom is array(0 to 4095) of std_logic_vector(7 downto 0);

signal rom : t_rom := (

-- Altair 4K Basic ROM as per file '4kbas32.bin' in the SIMH simulator

X"F3", X"C3", X"21", X"0D", X"90", X"04", X"F9", X"07", X"7E", X"E3", X"BE", X"23", X"E3", X"C2", X"D0", X"01",
X"23", X"7E", X"FE", X"3A", X"D0", X"C3", X"5E", X"04", X"F5", X"3A", X"27", X"00", X"C3", X"6E", X"03", X"00",
X"7C", X"92", X"C0", X"7D", X"93", X"C9", X"01", X"00", X"3A", X"72", X"01", X"B7", X"C2", X"DA", X"09", X"C9",
X"E3", X"22", X"3B", X"00", X"E1", X"4E", X"23", X"46", X"23", X"C5", X"C3", X"3A", X"00", X"E4", X"09", X"A2",
X"0A", X"F8", X"09", X"98", X"04", X"21", X"0C", X"5F", X"0C", X"95", X"0C", X"79", X"10", X"08", X"79", X"0A",
X"08", X"7C", X"E3", X"08", X"7C", X"2F", X"09", X"45", X"4E", X"C4", X"46", X"4F", X"D2", X"4E", X"45", X"58",
X"D4", X"44", X"41", X"54", X"C1", X"49", X"4E", X"50", X"55", X"D4", X"44", X"49", X"CD", X"52", X"45", X"41",
X"C4", X"4C", X"45", X"D4", X"47", X"4F", X"54", X"CF", X"52", X"55", X"CE", X"49", X"C6", X"52", X"45", X"53",
X"54", X"4F", X"52", X"C5", X"47", X"4F", X"53", X"55", X"C2", X"52", X"45", X"54", X"55", X"52", X"CE", X"52",
X"45", X"CD", X"53", X"54", X"4F", X"D0", X"50", X"52", X"49", X"4E", X"D4", X"4C", X"49", X"53", X"D4", X"43",
X"4C", X"45", X"41", X"D2", X"4E", X"45", X"D7", X"54", X"41", X"42", X"A8", X"54", X"CF", X"54", X"48", X"45",
X"CE", X"53", X"54", X"45", X"D0", X"AB", X"AD", X"AA", X"AF", X"BE", X"BD", X"BC", X"53", X"47", X"CE", X"49",
X"4E", X"D4", X"41", X"42", X"D3", X"55", X"53", X"D2", X"53", X"51", X"D2", X"52", X"4E", X"C4", X"53", X"49",
X"CE", X"00", X"F7", X"01", X"D5", X"03", X"49", X"06", X"F5", X"04", X"E4", X"05", X"16", X"07", X"F6", X"05",
X"02", X"05", X"CF", X"04", X"A1", X"02", X"16", X"05", X"69", X"04", X"BE", X"04", X"DF", X"04", X"F7", X"04",
X"F7", X"01", X"57", X"05", X"8E", X"03", X"A6", X"02", X"95", X"02", X"4E", X"C6", X"53", X"CE", X"52", X"C7",
X"4F", X"C4", X"46", X"C3", X"4F", X"D6", X"4F", X"CD", X"55", X"D3", X"42", X"D3", X"44", X"C4", X"2F", X"B0",
X"49", X"C4", X"2C", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"1A", X"0F", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"20", X"45", X"52", X"52", X"4F", X"D2", X"00", X"20", X"49", X"4E", X"A0", X"00", X"0D", X"4F", X"CB",
X"0D", X"00", X"21", X"04", X"00", X"39", X"7E", X"23", X"FE", X"81", X"C0", X"F7", X"E3", X"E7", X"01", X"0D",
X"00", X"E1", X"C8", X"09", X"C3", X"96", X"01", X"CD", X"C3", X"01", X"C5", X"E3", X"C1", X"E7", X"7E", X"02",
X"C8", X"0B", X"2B", X"C3", X"AD", X"01", X"E5", X"2A", X"6B", X"01", X"06", X"00", X"09", X"09", X"CD", X"C3",
X"01", X"E1", X"C9", X"D5", X"EB", X"21", X"DE", X"FF", X"39", X"E7", X"EB", X"D1", X"D0", X"1E", X"0C", X"01",
X"1E", X"02", X"01", X"1E", X"14", X"CD", X"B5", X"02", X"CD", X"8A", X"05", X"21", X"FA", X"00", X"57", X"3E",
X"3F", X"DF", X"19", X"7E", X"DF", X"D7", X"DF", X"21", X"81", X"01", X"CD", X"A3", X"05", X"2A", X"61", X"01",
X"7C", X"A5", X"3C", X"C4", X"2F", X"0B", X"01", X"C0", X"C1", X"21", X"8D", X"01", X"CD", X"21", X"0D", X"21",
X"FF", X"FF", X"22", X"61", X"01", X"CD", X"3C", X"03", X"D7", X"3C", X"3D", X"CA", X"FF", X"01", X"F5", X"CD",
X"9D", X"04", X"D5", X"CD", X"CC", X"02", X"47", X"D1", X"F1", X"D2", X"3E", X"04", X"D5", X"C5", X"D7", X"B7",
X"F5", X"CD", X"7D", X"02", X"C5", X"D2", X"39", X"02", X"EB", X"2A", X"67", X"01", X"1A", X"02", X"03", X"13",
X"E7", X"C2", X"2C", X"02", X"60", X"69", X"22", X"67", X"01", X"D1", X"F1", X"CA", X"60", X"02", X"2A", X"67",
X"01", X"E3", X"C1", X"09", X"E5", X"CD", X"A7", X"01", X"E1", X"22", X"67", X"01", X"EB", X"74", X"23", X"23",
X"D1", X"73", X"23", X"72", X"23", X"11", X"13", X"01", X"1A", X"77", X"23", X"13", X"B7", X"C2", X"58", X"02",
X"CD", X"A2", X"02", X"23", X"EB", X"62", X"6B", X"7E", X"23", X"B6", X"CA", X"FF", X"01", X"23", X"23", X"23",
X"AF", X"BE", X"23", X"C2", X"71", X"02", X"EB", X"73", X"23", X"72", X"C3", X"65", X"02", X"2A", X"65", X"01",
X"44", X"4D", X"7E", X"23", X"B6", X"2B", X"C8", X"C5", X"F7", X"F7", X"E1", X"E7", X"E1", X"C1", X"3F", X"C8",
X"3F", X"D0", X"C3", X"80", X"02", X"C0", X"2A", X"65", X"01", X"AF", X"77", X"23", X"77", X"23", X"22", X"67",
X"01", X"C0", X"2A", X"65", X"01", X"2B", X"22", X"5D", X"01", X"CD", X"69", X"04", X"2A", X"67", X"01", X"22",
X"69", X"01", X"22", X"6B", X"01", X"C1", X"2A", X"63", X"01", X"F9", X"AF", X"6F", X"E5", X"C5", X"2A", X"5D",
X"01", X"C9", X"3E", X"3F", X"DF", X"3E", X"20", X"DF", X"CD", X"3C", X"03", X"23", X"0E", X"05", X"11", X"13",
X"01", X"7E", X"FE", X"20", X"CA", X"02", X"03", X"47", X"FE", X"22", X"CA", X"15", X"03", X"B7", X"CA", X"29",
X"03", X"D5", X"06", X"00", X"11", X"56", X"00", X"E5", X"3E", X"D7", X"13", X"1A", X"E6", X"7F", X"CA", X"FF",
X"02", X"BE", X"C2", X"1C", X"03", X"1A", X"B7", X"F2", X"E9", X"02", X"F1", X"78", X"F6", X"80", X"F2", X"E1",
X"7E", X"D1", X"23", X"12", X"13", X"0C", X"D6", X"8E", X"C2", X"D1", X"02", X"47", X"7E", X"B7", X"CA", X"29",
X"03", X"B8", X"CA", X"02", X"03", X"23", X"12", X"0C", X"13", X"C3", X"0C", X"03", X"E1", X"E5", X"04", X"EB",
X"B6", X"23", X"F2", X"20", X"03", X"EB", X"C3", X"EB", X"02", X"21", X"12", X"01", X"12", X"13", X"12", X"13",
X"12", X"C9", X"05", X"2B", X"DF", X"C2", X"41", X"03", X"DF", X"CD", X"8A", X"05", X"21", X"13", X"01", X"06",
X"01", X"CD", X"82", X"03", X"FE", X"0D", X"CA", X"85", X"05", X"FE", X"20", X"DA", X"41", X"03", X"FE", X"7D",
X"D2", X"41", X"03", X"FE", X"40", X"CA", X"38", X"03", X"FE", X"5F", X"CA", X"32", X"03", X"4F", X"78", X"FE",
X"48", X"3E", X"07", X"D2", X"6A", X"03", X"79", X"71", X"23", X"04", X"DF", X"C3", X"41", X"03", X"FE", X"48",
X"CC", X"8A", X"05", X"3C", X"32", X"27", X"00", X"DB", X"00", X"E6", X"80", X"C2", X"77", X"03", X"F1", X"D3",
X"01", X"C9", X"DB", X"00", X"E6", X"01", X"C2", X"82", X"03", X"DB", X"01", X"E6", X"7F", X"C9", X"CD", X"9D",
X"04", X"C0", X"C1", X"CD", X"7D", X"02", X"C5", X"E1", X"F7", X"C1", X"78", X"B1", X"CA", X"F9", X"01", X"CD",
X"73", X"04", X"C5", X"CD", X"8A", X"05", X"F7", X"E3", X"CD", X"37", X"0B", X"3E", X"20", X"E1", X"DF", X"7E",
X"B7", X"23", X"CA", X"97", X"03", X"F2", X"AE", X"03", X"D6", X"7F", X"4F", X"E5", X"11", X"57", X"00", X"D5",
X"1A", X"13", X"B7", X"F2", X"C0", X"03", X"0D", X"E1", X"C2", X"BF", X"03", X"7E", X"B7", X"FA", X"AD", X"03",
X"DF", X"23", X"C3", X"CB", X"03", X"CD", X"02", X"05", X"E3", X"CD", X"92", X"01", X"D1", X"C2", X"E2", X"03",
X"09", X"F9", X"EB", X"0E", X"08", X"CD", X"B6", X"01", X"E5", X"CD", X"F5", X"04", X"E3", X"E5", X"2A", X"61",
X"01", X"E3", X"CF", X"95", X"CD", X"8A", X"06", X"E5", X"CD", X"1D", X"0A", X"E1", X"C5", X"D5", X"01", X"00",
X"81", X"51", X"5A", X"7E", X"FE", X"97", X"3E", X"01", X"C2", X"14", X"04", X"CD", X"8B", X"06", X"E5", X"CD",
X"1D", X"0A", X"EF", X"E1", X"C5", X"D5", X"F5", X"33", X"E5", X"2A", X"5D", X"01", X"E3", X"06", X"81", X"C5",
X"33", X"CD", X"73", X"04", X"7E", X"FE", X"3A", X"CA", X"3E", X"04", X"B7", X"C2", X"D0", X"01", X"23", X"7E",
X"23", X"B6", X"23", X"CA", X"F9", X"01", X"5E", X"23", X"56", X"EB", X"22", X"61", X"01", X"EB", X"D7", X"11",
X"21", X"04", X"D5", X"C8", X"D6", X"80", X"DA", X"02", X"05", X"FE", X"14", X"D2", X"D0", X"01", X"07", X"4F",
X"06", X"00", X"EB", X"21", X"D2", X"00", X"09", X"4E", X"23", X"46", X"C5", X"EB", X"D7", X"C9", X"FE", X"20",
X"CA", X"10", X"00", X"FE", X"30", X"3F", X"3C", X"3D", X"C9", X"EB", X"2A", X"65", X"01", X"2B", X"22", X"6D",
X"01", X"EB", X"C9", X"DB", X"00", X"E6", X"01", X"C0", X"CD", X"82", X"03", X"FE", X"03", X"C3", X"F7", X"01",
X"7E", X"FE", X"41", X"D8", X"FE", X"5B", X"3F", X"C9", X"D7", X"CD", X"8A", X"06", X"EF", X"FA", X"98", X"04",
X"3A", X"72", X"01", X"FE", X"90", X"DA", X"77", X"0A", X"1E", X"08", X"C3", X"D5", X"01", X"2B", X"11", X"00",
X"00", X"D7", X"D0", X"E5", X"F5", X"21", X"98", X"19", X"E7", X"DA", X"D0", X"01", X"62", X"6B", X"19", X"29",
X"19", X"29", X"F1", X"D6", X"30", X"5F", X"16", X"00", X"19", X"EB", X"E1", X"C3", X"A1", X"04", X"0E", X"03",
X"CD", X"B6", X"01", X"C1", X"E5", X"E5", X"2A", X"61", X"01", X"E3", X"16", X"8C", X"D5", X"33", X"C5", X"CD",
X"9D", X"04", X"C0", X"CD", X"7D", X"02", X"60", X"69", X"2B", X"D8", X"1E", X"0E", X"C3", X"D5", X"01", X"C0",
X"16", X"FF", X"CD", X"92", X"01", X"F9", X"FE", X"8C", X"1E", X"04", X"C2", X"D5", X"01", X"E1", X"22", X"61",
X"01", X"21", X"21", X"04", X"E3", X"01", X"3A", X"10", X"00", X"7E", X"B7", X"C8", X"B9", X"C8", X"23", X"C3",
X"F9", X"04", X"CD", X"1B", X"07", X"CF", X"9D", X"D5", X"CD", X"8A", X"06", X"E3", X"22", X"5D", X"01", X"E5",
X"CD", X"29", X"0A", X"D1", X"E1", X"C9", X"CD", X"8A", X"06", X"7E", X"CD", X"02", X"0A", X"16", X"00", X"D6",
X"9C", X"DA", X"32", X"05", X"FE", X"03", X"D2", X"32", X"05", X"FE", X"01", X"17", X"B2", X"57", X"D7", X"C3",
X"1F", X"05", X"7A", X"B7", X"CA", X"D0", X"01", X"F5", X"CD", X"8A", X"06", X"CF", X"96", X"2B", X"F1", X"C1",
X"D1", X"E5", X"F5", X"CD", X"4C", X"0A", X"3C", X"17", X"C1", X"A0", X"E1", X"CA", X"F7", X"04", X"D7", X"DA",
X"CF", X"04", X"C3", X"43", X"04", X"2B", X"D7", X"CA", X"8A", X"05", X"C8", X"FE", X"22", X"CC", X"A2", X"05",
X"CA", X"55", X"05", X"FE", X"94", X"CA", X"C7", X"05", X"E5", X"FE", X"2C", X"CA", X"B3", X"05", X"FE", X"3B",
X"CA", X"DF", X"05", X"C1", X"CD", X"8A", X"06", X"E5", X"CD", X"42", X"0B", X"CD", X"A3", X"05", X"3E", X"20",
X"DF", X"E1", X"C3", X"55", X"05", X"36", X"00", X"21", X"12", X"01", X"3E", X"0D", X"32", X"27", X"00", X"DF",
X"3E", X"0A", X"DF", X"3A", X"26", X"00", X"3D", X"32", X"27", X"00", X"C8", X"F5", X"AF", X"DF", X"F1", X"C3",
X"96", X"05", X"23", X"7E", X"B7", X"C8", X"23", X"FE", X"22", X"C8", X"DF", X"FE", X"0D", X"CC", X"8A", X"05",
X"C3", X"A3", X"05", X"3A", X"27", X"00", X"FE", X"38", X"D4", X"8A", X"05", X"D2", X"DF", X"05", X"D6", X"0E",
X"D2", X"BE", X"05", X"2F", X"C3", X"D6", X"05", X"CD", X"88", X"04", X"CF", X"29", X"2B", X"E5", X"3A", X"27",
X"00", X"2F", X"83", X"D2", X"DF", X"05", X"3C", X"47", X"3E", X"20", X"DF", X"05", X"C2", X"DA", X"05", X"E1",
X"D7", X"C3", X"5A", X"05", X"E5", X"2A", X"61", X"01", X"1E", X"16", X"23", X"7D", X"B4", X"CA", X"D5", X"01",
X"CD", X"C2", X"02", X"C3", X"FB", X"05", X"E5", X"2A", X"6D", X"01", X"F6", X"AF", X"32", X"5C", X"01", X"E3",
X"01", X"CF", X"2C", X"CD", X"1B", X"07", X"E3", X"D5", X"7E", X"FE", X"2C", X"CA", X"20", X"06", X"B7", X"C2",
X"D0", X"01", X"3A", X"5C", X"01", X"B7", X"23", X"C2", X"36", X"06", X"3E", X"3F", X"DF", X"CD", X"C2", X"02",
X"D1", X"23", X"CD", X"07", X"05", X"E3", X"2B", X"D7", X"C2", X"01", X"06", X"D1", X"3A", X"5C", X"01", X"B7",
X"C8", X"EB", X"C2", X"6E", X"04", X"E1", X"F7", X"79", X"B0", X"1E", X"06", X"CA", X"D5", X"01", X"23", X"D7",
X"FE", X"83", X"C2", X"35", X"06", X"C1", X"C3", X"20", X"06", X"CD", X"1B", X"07", X"22", X"5D", X"01", X"CD",
X"92", X"01", X"F9", X"D5", X"7E", X"23", X"F5", X"D5", X"1E", X"00", X"C2", X"D5", X"01", X"CD", X"0F", X"0A",
X"E3", X"E5", X"CD", X"04", X"08", X"E1", X"CD", X"29", X"0A", X"E1", X"CD", X"20", X"0A", X"E5", X"CD", X"4C",
X"0A", X"E1", X"C1", X"90", X"CD", X"20", X"0A", X"CA", X"83", X"06", X"EB", X"22", X"61", X"01", X"69", X"60",
X"C3", X"1D", X"04", X"F9", X"2A", X"5D", X"01", X"C3", X"21", X"04", X"2B", X"16", X"00", X"D5", X"0E", X"01",
X"CD", X"B6", X"01", X"CD", X"C4", X"06", X"22", X"5F", X"01", X"2A", X"5F", X"01", X"C1", X"7E", X"16", X"00",
X"D6", X"98", X"D8", X"FE", X"04", X"D0", X"5F", X"07", X"83", X"5F", X"21", X"4B", X"00", X"19", X"78", X"56",
X"BA", X"D0", X"23", X"C5", X"01", X"99", X"06", X"C5", X"4A", X"CD", X"02", X"0A", X"51", X"F7", X"2A", X"5F",
X"01", X"C3", X"8D", X"06", X"D7", X"DA", X"B3", X"0A", X"CD", X"80", X"04", X"D2", X"F3", X"06", X"FE", X"98",
X"CA", X"C4", X"06", X"FE", X"2E", X"CA", X"B3", X"0A", X"FE", X"99", X"CA", X"EA", X"06", X"D6", X"9F", X"D2",
X"FD", X"06", X"CF", X"28", X"CD", X"8A", X"06", X"CF", X"29", X"C9", X"CD", X"C4", X"06", X"E5", X"CD", X"FA",
X"09", X"E1", X"C9", X"CD", X"1B", X"07", X"E5", X"EB", X"CD", X"0F", X"0A", X"E1", X"C9", X"06", X"00", X"07",
X"4F", X"C5", X"D7", X"CD", X"E2", X"06", X"E3", X"11", X"F1", X"06", X"D5", X"01", X"3D", X"00", X"09", X"F7",
X"C9", X"2B", X"D7", X"C8", X"CF", X"2C", X"01", X"11", X"07", X"C5", X"F6", X"AF", X"32", X"5B", X"01", X"46",
X"CD", X"80", X"04", X"DA", X"D0", X"01", X"AF", X"4F", X"D7", X"D2", X"2E", X"07", X"4F", X"D7", X"D6", X"28",
X"CA", X"8A", X"07", X"E5", X"2A", X"69", X"01", X"EB", X"2A", X"67", X"01", X"E7", X"CA", X"52", X"07", X"79",
X"96", X"23", X"C2", X"47", X"07", X"78", X"96", X"23", X"CA", X"82", X"07", X"23", X"23", X"23", X"23", X"C3",
X"3B", X"07", X"E1", X"E3", X"D5", X"11", X"F6", X"06", X"E7", X"D1", X"CA", X"85", X"07", X"E3", X"E5", X"C5",
X"01", X"06", X"00", X"2A", X"6B", X"01", X"E5", X"09", X"C1", X"E5", X"CD", X"A7", X"01", X"E1", X"22", X"6B",
X"01", X"60", X"69", X"22", X"69", X"01", X"2B", X"36", X"00", X"E7", X"C2", X"76", X"07", X"D1", X"73", X"23",
X"72", X"23", X"EB", X"E1", X"C9", X"32", X"72", X"01", X"E1", X"C9", X"C5", X"3A", X"5B", X"01", X"F5", X"CD",
X"88", X"04", X"CF", X"29", X"F1", X"32", X"5B", X"01", X"E3", X"EB", X"29", X"29", X"E5", X"2A", X"69", X"01",
X"01", X"C1", X"09", X"EB", X"E5", X"2A", X"6B", X"01", X"E7", X"EB", X"D1", X"CA", X"CD", X"07", X"F7", X"E3",
X"E7", X"E1", X"F7", X"C2", X"A1", X"07", X"3A", X"5B", X"01", X"B7", X"1E", X"12", X"C2", X"D5", X"01", X"D1",
X"1B", X"E3", X"E7", X"1E", X"10", X"D2", X"D5", X"01", X"D1", X"19", X"D1", X"EB", X"C9", X"73", X"23", X"72",
X"23", X"11", X"2C", X"00", X"3A", X"5B", X"01", X"B7", X"CA", X"E1", X"07", X"D1", X"D5", X"13", X"13", X"13",
X"13", X"D5", X"73", X"23", X"72", X"23", X"E5", X"19", X"CD", X"C3", X"01", X"22", X"6B", X"01", X"D1", X"2B",
X"36", X"00", X"E7", X"C2", X"EF", X"07", X"C3", X"BF", X"07", X"50", X"1E", X"00", X"06", X"90", X"C3", X"EA",
X"09", X"21", X"0B", X"0C", X"CD", X"20", X"0A", X"C3", X"12", X"08", X"C1", X"D1", X"CD", X"FA", X"09", X"21",
X"C1", X"D1", X"78", X"B7", X"C8", X"3A", X"72", X"01", X"B7", X"CA", X"12", X"0A", X"90", X"D2", X"2C", X"08",
X"2F", X"3C", X"EB", X"CD", X"02", X"0A", X"EB", X"CD", X"12", X"0A", X"C1", X"D1", X"F5", X"CD", X"37", X"0A",
X"67", X"F1", X"CD", X"C9", X"08", X"B4", X"21", X"6F", X"01", X"F2", X"4D", X"08", X"CD", X"A9", X"08", X"D2",
X"7E", X"08", X"23", X"34", X"CA", X"A4", X"08", X"CD", X"D6", X"08", X"C3", X"7E", X"08", X"AF", X"90", X"47",
X"7E", X"9B", X"5F", X"23", X"7E", X"9A", X"57", X"23", X"7E", X"99", X"4F", X"DC", X"B5", X"08", X"26", X"00",
X"79", X"B7", X"FA", X"7E", X"08", X"FE", X"E0", X"CA", X"BE", X"09", X"25", X"78", X"87", X"47", X"CD", X"90",
X"08", X"7C", X"F2", X"65", X"08", X"21", X"72", X"01", X"86", X"77", X"D2", X"BE", X"09", X"C8", X"78", X"21",
X"72", X"01", X"B7", X"FC", X"9A", X"08", X"46", X"23", X"7E", X"E6", X"80", X"A9", X"4F", X"C3", X"12", X"0A",
X"7B", X"17", X"5F", X"7A", X"17", X"57", X"79", X"8F", X"4F", X"C9", X"1C", X"C0", X"14", X"C0", X"0C", X"C0",
X"0E", X"80", X"34", X"C0", X"1E", X"0A", X"C3", X"D5", X"01", X"7E", X"83", X"5F", X"23", X"7E", X"8A", X"57",
X"23", X"7E", X"89", X"4F", X"C9", X"21", X"73", X"01", X"7E", X"2F", X"77", X"AF", X"6F", X"90", X"47", X"7D",
X"9B", X"5F", X"7D", X"9A", X"57", X"7D", X"99", X"4F", X"C9", X"06", X"00", X"3C", X"6F", X"AF", X"2D", X"C8",
X"CD", X"D6", X"08", X"C3", X"CD", X"08", X"79", X"1F", X"4F", X"7A", X"1F", X"57", X"7B", X"1F", X"5F", X"78",
X"1F", X"47", X"C9", X"C1", X"D1", X"EF", X"C8", X"2E", X"00", X"CD", X"9B", X"09", X"79", X"32", X"17", X"09",
X"EB", X"22", X"12", X"09", X"01", X"00", X"00", X"50", X"58", X"21", X"5E", X"08", X"E5", X"21", X"05", X"09",
X"E5", X"E5", X"21", X"6F", X"01", X"7E", X"23", X"E5", X"2E", X"08", X"1F", X"67", X"79", X"D2", X"19", X"09",
X"E5", X"21", X"00", X"00", X"19", X"D1", X"CE", X"00", X"EB", X"CD", X"D7", X"08", X"2D", X"7C", X"C2", X"0A",
X"09", X"E1", X"C9", X"CD", X"02", X"0A", X"01", X"20", X"84", X"11", X"00", X"00", X"CD", X"12", X"0A", X"C1",
X"D1", X"EF", X"CA", X"D3", X"01", X"2E", X"FF", X"CD", X"9B", X"09", X"34", X"34", X"2B", X"7E", X"32", X"60",
X"09", X"2B", X"7E", X"32", X"5C", X"09", X"2B", X"7E", X"32", X"58", X"09", X"41", X"EB", X"AF", X"4F", X"57",
X"5F", X"32", X"63", X"09", X"E5", X"C5", X"7D", X"D6", X"00", X"6F", X"7C", X"DE", X"00", X"67", X"78", X"DE",
X"00", X"47", X"3E", X"00", X"DE", X"00", X"3F", X"D2", X"71", X"09", X"32", X"63", X"09", X"F1", X"F1", X"37",
X"D2", X"C1", X"E1", X"79", X"3C", X"3D", X"1F", X"FA", X"7F", X"08", X"17", X"CD", X"90", X"08", X"29", X"78",
X"17", X"47", X"3A", X"63", X"09", X"17", X"32", X"63", X"09", X"79", X"B2", X"B3", X"C2", X"54", X"09", X"E5",
X"21", X"72", X"01", X"35", X"E1", X"C2", X"54", X"09", X"C3", X"A4", X"08", X"78", X"B7", X"CA", X"BA", X"09",
X"7D", X"21", X"72", X"01", X"AE", X"80", X"47", X"1F", X"A8", X"78", X"F2", X"B9", X"09", X"C6", X"80", X"77",
X"CA", X"21", X"09", X"CD", X"37", X"0A", X"77", X"2B", X"C9", X"B7", X"E1", X"FA", X"A4", X"08", X"AF", X"32",
X"72", X"01", X"C9", X"CD", X"1D", X"0A", X"78", X"B7", X"C8", X"C6", X"02", X"DA", X"A4", X"08", X"47", X"CD",
X"12", X"08", X"21", X"72", X"01", X"34", X"C0", X"C3", X"A4", X"08", X"3A", X"71", X"01", X"FE", X"2F", X"17",
X"9F", X"C0", X"3C", X"C9", X"EF", X"06", X"88", X"11", X"00", X"00", X"21", X"72", X"01", X"4F", X"70", X"06",
X"00", X"23", X"36", X"80", X"17", X"C3", X"5B", X"08", X"EF", X"F0", X"21", X"71", X"01", X"7E", X"EE", X"80",
X"77", X"C9", X"EB", X"2A", X"6F", X"01", X"E3", X"E5", X"2A", X"71", X"01", X"E3", X"E5", X"EB", X"C9", X"CD",
X"20", X"0A", X"EB", X"22", X"6F", X"01", X"60", X"69", X"22", X"71", X"01", X"EB", X"C9", X"21", X"6F", X"01",
X"5E", X"23", X"56", X"23", X"4E", X"23", X"46", X"23", X"C9", X"11", X"6F", X"01", X"06", X"04", X"1A", X"77",
X"13", X"23", X"05", X"C2", X"2E", X"0A", X"C9", X"21", X"71", X"01", X"7E", X"07", X"37", X"1F", X"77", X"3F",
X"1F", X"23", X"23", X"77", X"79", X"07", X"37", X"1F", X"4F", X"1F", X"AE", X"C9", X"78", X"B7", X"CA", X"28",
X"00", X"21", X"DE", X"09", X"E5", X"EF", X"79", X"C8", X"21", X"71", X"01", X"AE", X"79", X"F8", X"CD", X"64",
X"0A", X"1F", X"A9", X"C9", X"23", X"78", X"BE", X"C0", X"2B", X"79", X"BE", X"C0", X"2B", X"7A", X"BE", X"C0",
X"2B", X"7B", X"96", X"C0", X"E1", X"E1", X"C9", X"47", X"4F", X"57", X"5F", X"B7", X"C8", X"E5", X"CD", X"1D",
X"0A", X"CD", X"37", X"0A", X"AE", X"67", X"FC", X"9B", X"0A", X"3E", X"98", X"90", X"CD", X"C9", X"08", X"7C",
X"17", X"DC", X"9A", X"08", X"06", X"00", X"DC", X"B5", X"08", X"E1", X"C9", X"1B", X"7A", X"A3", X"3C", X"C0",
X"0D", X"C9", X"21", X"72", X"01", X"7E", X"FE", X"98", X"D0", X"CD", X"77", X"0A", X"36", X"98", X"79", X"17",
X"C3", X"5B", X"08", X"2B", X"CD", X"BE", X"09", X"47", X"57", X"5F", X"2F", X"4F", X"D7", X"DA", X"04", X"0B",
X"FE", X"2E", X"CA", X"E4", X"0A", X"FE", X"45", X"C2", X"E8", X"0A", X"D7", X"15", X"FE", X"99", X"CA", X"D8",
X"0A", X"14", X"FE", X"98", X"CA", X"D8", X"0A", X"2B", X"D7", X"DA", X"23", X"0B", X"14", X"C2", X"E8", X"0A",
X"AF", X"93", X"5F", X"0C", X"0C", X"CA", X"BC", X"0A", X"E5", X"7B", X"90", X"F4", X"FC", X"0A", X"F2", X"F7",
X"0A", X"F5", X"CD", X"23", X"09", X"F1", X"3C", X"C2", X"EB", X"0A", X"E1", X"C9", X"C8", X"F5", X"CD", X"C3",
X"09", X"F1", X"3D", X"C9", X"D5", X"57", X"78", X"89", X"47", X"C5", X"E5", X"D5", X"CD", X"C3", X"09", X"F1",
X"D6", X"30", X"CD", X"02", X"0A", X"CD", X"E5", X"09", X"C1", X"D1", X"CD", X"12", X"08", X"E1", X"C1", X"D1",
X"C3", X"BC", X"0A", X"7B", X"07", X"07", X"83", X"07", X"86", X"D6", X"30", X"5F", X"C3", X"D8", X"0A", X"E5",
X"21", X"88", X"01", X"CD", X"A3", X"05", X"E1", X"EB", X"AF", X"06", X"98", X"CD", X"EA", X"09", X"21", X"A2",
X"05", X"E5", X"21", X"74", X"01", X"E5", X"EF", X"36", X"20", X"F2", X"4E", X"0B", X"36", X"2D", X"23", X"36",
X"30", X"CA", X"F7", X"0B", X"E5", X"FC", X"FA", X"09", X"AF", X"F5", X"CD", X"FD", X"0B", X"01", X"43", X"91",
X"11", X"F8", X"4F", X"CD", X"4C", X"0A", X"E2", X"7A", X"0B", X"F1", X"CD", X"FD", X"0A", X"F5", X"C3", X"5D",
X"0B", X"CD", X"23", X"09", X"F1", X"3C", X"F5", X"CD", X"FD", X"0B", X"CD", X"01", X"08", X"3C", X"CD", X"77",
X"0A", X"CD", X"12", X"0A", X"01", X"06", X"02", X"F1", X"81", X"FA", X"95", X"0B", X"FE", X"07", X"D2", X"95",
X"0B", X"3C", X"47", X"3E", X"01", X"3D", X"E1", X"F5", X"11", X"0F", X"0C", X"05", X"36", X"2E", X"CC", X"27",
X"0A", X"C5", X"E5", X"D5", X"CD", X"1D", X"0A", X"E1", X"06", X"2F", X"04", X"7B", X"96", X"5F", X"23", X"7A",
X"9E", X"57", X"23", X"79", X"9E", X"4F", X"2B", X"2B", X"D2", X"AA", X"0B", X"CD", X"A9", X"08", X"23", X"CD",
X"12", X"0A", X"EB", X"E1", X"70", X"23", X"C1", X"0D", X"C2", X"9B", X"0B", X"05", X"CA", X"DB", X"0B", X"2B",
X"7E", X"FE", X"30", X"CA", X"CF", X"0B", X"FE", X"2E", X"C4", X"27", X"0A", X"F1", X"CA", X"FA", X"0B", X"36",
X"45", X"23", X"36", X"2B", X"F2", X"EB", X"0B", X"36", X"2D", X"2F", X"3C", X"06", X"2F", X"04", X"D6", X"0A",
X"D2", X"ED", X"0B", X"C6", X"3A", X"23", X"70", X"23", X"77", X"23", X"71", X"E1", X"C9", X"01", X"74", X"94",
X"11", X"F7", X"23", X"CD", X"4C", X"0A", X"E1", X"E2", X"71", X"0B", X"E9", X"00", X"00", X"00", X"80", X"A0",
X"86", X"01", X"10", X"27", X"00", X"E8", X"03", X"00", X"64", X"00", X"00", X"0A", X"00", X"00", X"01", X"00",
X"00", X"EF", X"FA", X"98", X"04", X"C8", X"21", X"72", X"01", X"7E", X"1F", X"F5", X"E5", X"3E", X"40", X"17",
X"77", X"21", X"74", X"01", X"CD", X"29", X"0A", X"3E", X"04", X"F5", X"CD", X"02", X"0A", X"21", X"74", X"01",
X"CD", X"20", X"0A", X"CD", X"31", X"09", X"C1", X"D1", X"CD", X"12", X"08", X"01", X"00", X"80", X"51", X"59",
X"CD", X"E5", X"08", X"F1", X"3D", X"C2", X"39", X"0C", X"E1", X"F1", X"C6", X"C0", X"86", X"77", X"C9", X"EF",
X"FA", X"7C", X"0C", X"21", X"91", X"0C", X"CD", X"0F", X"0A", X"C8", X"01", X"35", X"98", X"11", X"7A", X"44",
X"CD", X"E5", X"08", X"01", X"28", X"68", X"11", X"46", X"B1", X"CD", X"12", X"08", X"CD", X"1D", X"0A", X"7B",
X"59", X"4F", X"36", X"80", X"2B", X"46", X"36", X"80", X"CD", X"5E", X"08", X"21", X"91", X"0C", X"C3", X"29",
X"0A", X"52", X"C7", X"4F", X"80", X"CD", X"02", X"0A", X"01", X"49", X"83", X"11", X"DB", X"0F", X"CD", X"12",
X"0A", X"C1", X"D1", X"CD", X"31", X"09", X"CD", X"02", X"0A", X"CD", X"A2", X"0A", X"C1", X"D1", X"CD", X"0C",
X"08", X"01", X"00", X"7F", X"51", X"59", X"CD", X"0C", X"08", X"EF", X"37", X"F2", X"C3", X"0C", X"CD", X"01",
X"08", X"EF", X"B7", X"F5", X"F4", X"FA", X"09", X"01", X"00", X"7F", X"51", X"59", X"CD", X"12", X"08", X"F1",
X"D4", X"FA", X"09", X"CD", X"02", X"0A", X"CD", X"1D", X"0A", X"CD", X"E5", X"08", X"CD", X"02", X"0A", X"21",
X"03", X"0D", X"CD", X"0F", X"0A", X"C1", X"D1", X"3E", X"04", X"F5", X"D5", X"C5", X"E5", X"CD", X"E5", X"08",
X"E1", X"CD", X"20", X"0A", X"E5", X"CD", X"12", X"08", X"E1", X"C1", X"D1", X"F1", X"3D", X"C2", X"E9", X"0C",
X"C3", X"E3", X"08", X"BA", X"D7", X"1E", X"86", X"64", X"26", X"99", X"87", X"58", X"34", X"23", X"87", X"E0",
X"5D", X"A5", X"86", X"DA", X"0F", X"49", X"83", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"21", X"1A", X"0F", X"F9", X"22", X"63", X"01", X"DB", X"01", X"0E", X"FF", X"11", X"8E", X"0D", X"D5",
X"3A", X"FF", X"0F", X"47", X"DB", X"FF", X"1F", X"DA", X"41", X"0D", X"E6", X"0C", X"CA", X"42", X"0D", X"06",
X"10", X"78", X"32", X"8C", X"0D", X"DB", X"FF", X"17", X"17", X"06", X"20", X"11", X"02", X"CA", X"D8", X"17",
X"43", X"1D", X"D8", X"17", X"DA", X"6F", X"0D", X"43", X"11", X"80", X"C2", X"17", X"D0", X"17", X"3E", X"03",
X"CD", X"8B", X"0D", X"3D", X"8F", X"87", X"87", X"3C", X"CD", X"8B", X"0D", X"37", X"C3", X"4B", X"0D", X"AF",
X"CD", X"8B", X"0D", X"CD", X"87", X"0D", X"CD", X"87", X"0D", X"4B", X"2F", X"CD", X"87", X"0D", X"3E", X"04",
X"35", X"CD", X"8B", X"0D", X"35", X"35", X"35", X"21", X"8C", X"0D", X"34", X"D3", X"10", X"C9", X"62", X"68",
X"22", X"85", X"03", X"7C", X"E6", X"C8", X"67", X"22", X"76", X"04", X"EB", X"22", X"7A", X"03", X"3A", X"8C",
X"0D", X"32", X"83", X"03", X"32", X"74", X"04", X"3C", X"32", X"8A", X"03", X"81", X"32", X"78", X"03", X"3C",
X"32", X"80", X"03", X"21", X"FF", X"FF", X"22", X"61", X"01", X"CD", X"8A", X"05", X"21", X"F0", X"0E", X"CD",
X"A3", X"05", X"CD", X"C2", X"02", X"D7", X"B7", X"C2", X"DE", X"0D", X"21", X"FC", X"0E", X"23", X"3E", X"37",
X"77", X"BE", X"C2", X"EA", X"0D", X"3D", X"77", X"BE", X"CA", X"CD", X"0D", X"C3", X"EA", X"0D", X"21", X"13",
X"01", X"CD", X"9D", X"04", X"B7", X"C2", X"D0", X"01", X"EB", X"2B", X"2B", X"E5", X"21", X"B4", X"0E", X"CD",
X"A3", X"05", X"CD", X"C2", X"02", X"D7", X"B7", X"CA", X"1B", X"0E", X"21", X"13", X"01", X"CD", X"9D", X"04",
X"7A", X"B7", X"C2", X"EC", X"0D", X"7B", X"FE", X"10", X"DA", X"EC", X"0D", X"32", X"6F", X"03", X"D6", X"0E",
X"D2", X"0E", X"0E", X"C6", X"1C", X"2F", X"3C", X"83", X"32", X"B7", X"05", X"21", X"85", X"0E", X"F7", X"11",
X"99", X"0E", X"E7", X"CA", X"32", X"0E", X"F7", X"E3", X"CD", X"A3", X"05", X"CD", X"C2", X"02", X"D7", X"E1",
X"FE", X"59", X"D1", X"CA", X"47", X"0E", X"FE", X"4E", X"C2", X"1B", X"0E", X"F7", X"E3", X"11", X"98", X"04",
X"73", X"23", X"72", X"E1", X"C3", X"1E", X"0E", X"EB", X"36", X"00", X"23", X"22", X"65", X"01", X"E3", X"11",
X"1A", X"0F", X"E7", X"DA", X"CD", X"01", X"D1", X"F9", X"22", X"63", X"01", X"EB", X"CD", X"C3", X"01", X"7B",
X"95", X"6F", X"7A", X"9C", X"67", X"01", X"F0", X"FF", X"09", X"CD", X"8A", X"05", X"CD", X"37", X"0B", X"21",
X"C3", X"0E", X"CD", X"A3", X"05", X"21", X"A3", X"05", X"22", X"FD", X"01", X"CD", X"96", X"02", X"21", X"F9",
X"01", X"22", X"02", X"00", X"E9", X"17", X"0D", X"99", X"0E", X"49", X"00", X"95", X"0C", X"A2", X"0E", X"47",
X"00", X"5F", X"0C", X"AB", X"0E", X"45", X"00", X"21", X"0C", X"57", X"41", X"4E", X"54", X"20", X"53", X"49",
X"CE", X"00", X"57", X"41", X"4E", X"54", X"20", X"52", X"4E", X"C4", X"00", X"57", X"41", X"4E", X"54", X"20",
X"53", X"51", X"D2", X"00", X"54", X"45", X"52", X"4D", X"49", X"4E", X"41", X"4C", X"20", X"57", X"49", X"44",
X"54", X"C8", X"00", X"20", X"42", X"59", X"54", X"45", X"53", X"20", X"46", X"52", X"45", X"C5", X"0D", X"0D",
X"42", X"41", X"53", X"49", X"43", X"20", X"56", X"45", X"52", X"53", X"49", X"4F", X"4E", X"20", X"33", X"2E",
X"B2", X"0D", X"5B", X"34", X"4B", X"20", X"56", X"45", X"52", X"53", X"49", X"4F", X"4E", X"DD", X"0D", X"00",
X"4D", X"45", X"4D", X"4F", X"52", X"59", X"20", X"53", X"49", X"5A", X"C5", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"

);


begin


rom_addr <= addr(11 downto 0);
process(clk)
begin
  if (clk'event and clk='1') then
    if we='1' then
      rom(conv_integer(rom_addr)) <= data_in;
    end if;
    data_out <= rom(conv_integer(rom_addr));
  end if;
end process;

end internal;
