/*
Developed By Subtleware Corporation Pte Ltd 2011
File		:
Description	:	
Remarks		:
Revision	:
	Date	Author		Description
02/09/12	Jefflieu
*/

module mClkBuf(input i_Clk,output o_Clk);

	
	assign o_Clk = i_Clk;
endmodule
