// megafunction wizard: %FIFO%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: scfifo

// ============================================================
// File Name: sc_fifo.v
// Megafunction Name(s):
// 			scfifo
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 7.2 Build 175 11/20/2007 SP 1 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2007 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions
//and other software and tools, and its AMPP partner logic
//functions, and any output files from any of the foregoing
//(including device programming or simulation files), and any
//associated documentation or information are expressly subject
//to the terms and conditions of the Altera Program License
//Subscription Agreement, Altera MegaCore Function License
//Agreement, or other applicable license agreement, including,
//without limitation, that your use is for the sole purpose of
//programming logic devices manufactured by Altera and sold by
//Altera or its authorized distributors.  Please refer to the
//applicable agreement for further details.

module alt_scfifo (
   aclr,
   clock,
   data,
   rdreq,
   sclr,
   wrreq,
   almost_empty,
   almost_full,
   empty,
   full,
   q,
   usedw,
   fifo_ovf,
   fifo_unf
);

   parameter                 FIFO_WIDTH    = 144;
   parameter                 FIFO_DEPTH    = 7;
   parameter                 FIFO_TYPE     = "AUTO";
   parameter                 FIFO_SHOW     = "OFF";
   parameter                 USE_EAB       = "ON";

   parameter                 FIFO_NUMWORDS = 1 << FIFO_DEPTH;
   parameter                 FIFO_AEMPTY   = 0;
   parameter                 FIFO_AFULL    = FIFO_NUMWORDS;
   parameter                 FIFO_UNF      = "TRUE";

   parameter                 TYPE          = FIFO_TYPE == "M4K"   | FIFO_TYPE == "M9K"  ?  "RAM_BLOCK_TYPE=M9K":
                                             FIFO_TYPE == "M512"  | FIFO_TYPE == "MLAB" ?  "RAM_BLOCK_TYPE=MLAB":
                                             FIFO_TYPE == "M-RAM" | FIFO_TYPE == "M144K"?  "RAM_BLOCK_TYPE=M144K":
                                                                                           "RAM_BLOCK_TYPE=AUTO";

   input                     aclr;
   input                     clock;
   input [FIFO_WIDTH-1:0]    data;
   input                     rdreq;
   input                     sclr;
   input                     wrreq;
   output                    almost_empty;
   output                    almost_full;
   output                    empty;
   output                    full;
   output [FIFO_WIDTH-1:0]   q;
   output [FIFO_DEPTH-1:0]   usedw;
   output                    fifo_ovf;
   output                    fifo_unf;

   reg                       fifo_ovf;
   reg                       fifo_unf;

   always @ (posedge clock or posedge aclr)
     if (aclr) begin
        fifo_ovf <= 1'b0;
        fifo_unf <= 1'b0;
     end
     else begin
        // synthesis translate_off
        if (fifo_ovf) begin
           $display ("%m: ERROR!!! %m alt_scfifo FIFO overflow, simulation stop");
           $stop;
        end
        if (fifo_unf & (FIFO_UNF == "TRUE")) begin
           $display ("%m: ERROR!!! alt_dcfifo FIFO underflow, simulation stop");
           $stop;
        end
        // synthesis translate_on
        fifo_ovf <=  (full  & wrreq) | fifo_ovf;
        fifo_unf <= ((empty & rdreq) | fifo_unf) & (FIFO_UNF == "TRUE");
     end

   scfifo scfifo_component (
      .rdreq       (rdreq),
      .sclr        (sclr),
      .aclr        (aclr),
      .clock       (clock),
      .wrreq       (wrreq),
      .data        (data),
      .almost_full (almost_full),
      .usedw       (usedw),
      .empty       (empty),
      .almost_empty(almost_empty),
      .q           (q),
      .full        (full)
      );
   defparam
	   scfifo_component.add_ram_output_register = "ON",
	   scfifo_component.almost_empty_value = FIFO_AEMPTY,
	   scfifo_component.almost_full_value = FIFO_AFULL,
	   scfifo_component.intended_device_family = "Stratix III",
	   scfifo_component.lpm_hint = TYPE,
	   scfifo_component.lpm_numwords = FIFO_NUMWORDS,
	   scfifo_component.lpm_showahead = FIFO_SHOW,
	   scfifo_component.lpm_type = "scfifo",
	   scfifo_component.lpm_width = FIFO_WIDTH,
	   scfifo_component.lpm_widthu = FIFO_DEPTH,
	   scfifo_component.overflow_checking = "ON",
	   scfifo_component.underflow_checking = "ON",
	   scfifo_component.use_eab = USE_EAB;
endmodule // alt_scfifo
