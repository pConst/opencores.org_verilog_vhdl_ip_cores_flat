-- obj_code_pkg -- Object code in VHDL constant table for BRAM initialization.
-- Generated automatically with script 'build_rom.py'.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.l80pkg.all;

package obj_code_pkg is

constant obj_code : obj_code_t(0 to 4848) := (
    X"c3", X"00", X"01", X"00", X"00", X"c3", X"a6", X"0e", 
    X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c3", X"13", X"01", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"21", X"40", X"1f", X"f9", X"11", 
    X"f8", X"0d", X"0e", X"09", X"cd", X"ec", X"0d", X"21", 
    X"3c", X"01", X"7e", X"23", X"b6", X"ca", X"2f", X"01", 
    X"2b", X"cd", X"d0", X"0a", X"c3", X"22", X"01", X"11", 
    X"15", X"0e", X"0e", X"09", X"cd", X"ec", X"0d", X"f3", 
    X"76", X"c3", X"00", X"00", X"70", X"01", X"d0", X"01", 
    X"30", X"02", X"90", X"02", X"f0", X"02", X"50", X"03", 
    X"b0", X"03", X"10", X"04", X"70", X"04", X"d0", X"04", 
    X"30", X"05", X"90", X"05", X"f0", X"05", X"50", X"06", 
    X"b0", X"06", X"10", X"07", X"70", X"07", X"d0", X"07", 
    X"30", X"08", X"90", X"08", X"f0", X"08", X"50", X"09", 
    X"b0", X"09", X"10", X"0a", X"70", X"0a", X"00", X"00", 
    X"ff", X"09", X"00", X"00", X"00", X"a5", X"c4", X"c7", 
    X"c4", X"26", X"d2", X"50", X"a0", X"ea", X"58", X"66", 
    X"85", X"c6", X"de", X"c9", X"9b", X"30", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"21", 
    X"f8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"ff", X"ff", X"ff", X"ff", X"ff", 
    X"ff", X"d7", X"00", X"ff", X"ff", X"14", X"47", X"4b", 
    X"a6", X"64", X"61", X"64", X"20", X"3c", X"62", X"2c", 
    X"64", X"2c", X"68", X"2c", X"73", X"70", X"3e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"c6", X"00", X"00", X"00", X"40", X"91", X"3c", 
    X"7e", X"67", X"7a", X"6d", X"df", X"61", X"5b", X"29", 
    X"0b", X"10", X"66", X"b2", X"85", X"38", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"ff", X"00", 
    X"00", X"00", X"ff", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"9e", X"92", X"2f", 
    X"9e", X"61", X"6c", X"75", X"6f", X"70", X"20", X"6e", 
    X"6e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"80", X"00", X"00", X"00", X"3e", X"c5", X"3a", 
    X"57", X"4d", X"4c", X"03", X"01", X"09", X"e3", X"66", 
    X"a6", X"d0", X"3b", X"bb", X"ad", X"3f", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"ff", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"ff", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"ff", X"ff", X"ff", 
    X"ff", X"d7", X"00", X"00", X"00", X"cf", X"76", X"2c", 
    X"86", X"61", X"6c", X"75", X"6f", X"70", X"20", X"3c", 
    X"62", X"2c", X"63", X"2c", X"64", X"2c", X"65", X"2c", 
    X"68", X"2c", X"6c", X"2c", X"6d", X"2c", X"61", X"3e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"27", X"00", X"00", X"00", X"41", X"21", X"fa", 
    X"09", X"60", X"1d", X"59", X"a5", X"5b", X"8d", X"79", 
    X"90", X"04", X"8e", X"9d", X"29", X"18", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"d7", X"ff", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"bb", X"3f", X"03", 
    X"0c", X"3c", X"64", X"61", X"61", X"2c", X"63", X"6d", 
    X"61", X"2c", X"73", X"74", X"63", X"2c", X"63", X"6d", 
    X"63", X"3e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"3c", X"00", X"00", X"00", X"df", X"4a", X"d8", 
    X"d5", X"98", X"e5", X"2b", X"8a", X"b0", X"a7", X"1b", 
    X"43", X"44", X"5a", X"30", X"d0", X"01", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"ff", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"ad", X"b6", X"46", 
    X"0e", X"3c", X"69", X"6e", X"72", X"2c", X"64", X"63", 
    X"72", X"3e", X"20", X"61", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"04", X"00", X"00", X"00", X"23", X"d6", X"2d", 
    X"43", X"61", X"7a", X"80", X"81", X"86", X"5a", X"85", 
    X"1e", X"86", X"58", X"bb", X"9b", X"01", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"ff", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"83", X"ed", X"13", 
    X"45", X"3c", X"69", X"6e", X"72", X"2c", X"64", X"63", 
    X"72", X"3e", X"20", X"62", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"03", X"00", X"00", X"00", X"97", X"cd", X"ab", 
    X"44", X"c9", X"8d", X"e3", X"e3", X"cc", X"11", X"a4", 
    X"e8", X"02", X"49", X"4d", X"2a", X"08", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"21", X"f8", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"f7", X"92", X"87", 
    X"cd", X"3c", X"69", X"6e", X"78", X"2c", X"64", X"63", 
    X"78", X"3e", X"20", X"62", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"0c", X"00", X"00", X"00", X"89", X"d7", X"35", 
    X"09", X"5b", X"05", X"85", X"9f", X"27", X"8b", X"08", 
    X"d2", X"95", X"05", X"60", X"06", X"01", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"ff", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"e5", X"f6", X"72", 
    X"1b", X"3c", X"69", X"6e", X"72", X"2c", X"64", X"63", 
    X"72", X"3e", X"20", X"63", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"14", X"00", X"00", X"00", X"ea", X"a0", X"ba", 
    X"5f", X"fb", X"65", X"1c", X"98", X"cc", X"38", X"bc", 
    X"de", X"43", X"5c", X"bd", X"03", X"01", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"ff", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"15", X"b5", X"57", 
    X"9a", X"3c", X"69", X"6e", X"72", X"2c", X"64", X"63", 
    X"72", X"3e", X"20", X"64", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"13", X"00", X"00", X"00", X"2e", X"34", X"1d", 
    X"13", X"c9", X"28", X"ca", X"0a", X"67", X"99", X"2e", 
    X"3a", X"92", X"f6", X"54", X"9d", X"08", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"21", X"f8", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"7f", X"4e", X"25", 
    X"01", X"3c", X"69", X"6e", X"78", X"2c", X"64", X"63", 
    X"78", X"3e", X"20", X"64", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"1c", X"00", X"00", X"00", X"2f", X"60", X"0d", 
    X"4c", X"02", X"24", X"f5", X"e2", X"f4", X"a0", X"0a", 
    X"a1", X"13", X"32", X"25", X"59", X"01", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"ff", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"cf", X"2a", X"b3", 
    X"96", X"3c", X"69", X"6e", X"72", X"2c", X"64", X"63", 
    X"72", X"3e", X"20", X"65", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"24", X"00", X"00", X"00", X"06", X"15", X"eb", 
    X"f2", X"dd", X"e8", X"2b", X"26", X"a6", X"11", X"1a", 
    X"bc", X"17", X"06", X"18", X"28", X"01", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"ff", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"12", X"b2", X"95", 
    X"2c", X"3c", X"69", X"6e", X"72", X"2c", X"64", X"63", 
    X"72", X"3e", X"20", X"68", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"23", X"00", X"00", X"00", X"f4", X"c3", X"a5", 
    X"07", X"6d", X"1b", X"04", X"4f", X"c2", X"e2", X"2a", 
    X"82", X"57", X"e0", X"e1", X"c3", X"08", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"21", 
    X"f8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"9f", X"2b", X"23", 
    X"c0", X"3c", X"69", X"6e", X"78", X"2c", X"64", X"63", 
    X"78", X"3e", X"20", X"68", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"2c", X"00", X"00", X"00", X"31", X"80", X"20", 
    X"a5", X"56", X"43", X"09", X"b4", X"c1", X"f4", X"a2", 
    X"df", X"d1", X"3c", X"a2", X"3e", X"01", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"ff", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"ff", X"57", X"d3", 
    X"56", X"3c", X"69", X"6e", X"72", X"2c", X"64", X"63", 
    X"72", X"3e", X"20", X"6c", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"34", X"00", X"00", X"00", X"56", X"b8", X"7c", 
    X"0c", X"3e", X"e5", X"03", X"01", X"7e", X"87", X"58", 
    X"da", X"15", X"5c", X"37", X"1f", X"01", X"00", X"00", 
    X"00", X"ff", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"92", X"e9", X"63", 
    X"bd", X"3c", X"69", X"6e", X"72", X"2c", X"64", X"63", 
    X"72", X"3e", X"20", X"6d", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"33", X"00", X"00", X"00", X"6f", X"34", X"82", 
    X"d4", X"69", X"d1", X"b6", X"de", X"94", X"a4", X"76", 
    X"f4", X"53", X"02", X"5b", X"85", X"08", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"21", 
    X"f8", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"d5", X"70", X"2f", 
    X"ab", X"3c", X"69", X"6e", X"78", X"2c", X"64", X"63", 
    X"78", X"3e", X"20", X"73", X"70", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"2a", X"03", X"01", X"00", X"63", X"98", X"30", 
    X"78", X"77", X"20", X"fe", X"b1", X"fa", X"b9", X"b8", 
    X"ab", X"04", X"06", X"15", X"60", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"ff", X"ff", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"a9", X"c3", X"d5", 
    X"cb", X"6c", X"68", X"6c", X"64", X"20", X"6e", X"6e", 
    X"6e", X"6e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"22", X"03", X"01", X"00", X"03", X"d0", X"72", 
    X"77", X"53", X"7f", X"72", X"3f", X"ea", X"64", X"80", 
    X"e1", X"10", X"2d", X"e9", X"35", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"ff", X"ff", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"e8", X"86", X"4f", 
    X"26", X"73", X"68", X"6c", X"64", X"20", X"6e", X"6e", 
    X"6e", X"6e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"01", X"00", X"00", X"00", X"1c", X"5c", X"46", 
    X"2d", X"b9", X"8e", X"78", X"60", X"b1", X"74", X"0e", 
    X"b3", X"46", X"d1", X"cc", X"30", X"30", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"ff", X"ff", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"fc", X"f4", X"6e", 
    X"12", X"6c", X"78", X"69", X"20", X"3c", X"62", X"2c", 
    X"64", X"2c", X"68", X"2c", X"73", X"70", X"3e", X"2c", 
    X"6e", X"6e", X"6e", X"6e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"0a", X"00", X"00", X"00", X"a8", X"b3", X"2a", 
    X"1d", X"8e", X"7f", X"ac", X"42", X"03", X"01", X"03", 
    X"01", X"c6", X"b1", X"8e", X"ef", X"10", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"ff", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"ff", X"00", X"00", X"2b", X"82", X"1d", 
    X"5f", X"6c", X"64", X"61", X"78", X"20", X"3c", X"62", 
    X"2c", X"64", X"3e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"06", X"00", X"00", X"00", X"07", X"c4", X"9d", 
    X"f4", X"3d", X"d1", X"39", X"03", X"89", X"de", X"55", 
    X"74", X"53", X"c0", X"09", X"55", X"38", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"ff", X"00", X"00", X"ea", X"a7", X"20", 
    X"44", X"6d", X"76", X"69", X"20", X"3c", X"62", X"2c", 
    X"63", X"2c", X"64", X"2c", X"65", X"2c", X"68", X"2c", 
    X"6c", X"2c", X"6d", X"2c", X"61", X"3e", X"2c", X"6e", 
    X"6e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"40", X"00", X"00", X"00", X"a4", X"72", X"24", 
    X"a0", X"ac", X"61", X"03", X"01", X"c7", X"82", X"8f", 
    X"71", X"97", X"8f", X"8e", X"ef", X"3f", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"ff", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"ff", X"ff", X"ff", 
    X"ff", X"d7", X"ff", X"00", X"00", X"10", X"b5", X"8c", 
    X"ee", X"6d", X"6f", X"76", X"20", X"3c", X"62", X"63", 
    X"64", X"65", X"68", X"6c", X"61", X"3e", X"2c", X"3c", 
    X"62", X"63", X"64", X"65", X"68", X"6c", X"61", X"3e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"32", X"03", X"01", X"00", X"68", X"fd", X"ec", 
    X"f4", X"a0", X"44", X"43", X"b5", X"53", X"06", X"ba", 
    X"cd", X"d2", X"4f", X"d8", X"1f", X"08", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"ff", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"ff", X"00", X"00", X"ed", X"57", X"af", 
    X"72", X"73", X"74", X"61", X"20", X"6e", X"6e", X"6e", 
    X"6e", X"20", X"2f", X"20", X"6c", X"64", X"61", X"20", 
    X"6e", X"6e", X"6e", X"6e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"07", X"00", X"00", X"00", X"92", X"cb", X"43", 
    X"6d", X"90", X"0a", X"84", X"c2", X"53", X"0c", X"0e", 
    X"f5", X"91", X"eb", X"fc", X"40", X"18", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"ff", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"d7", X"00", X"00", X"00", X"e0", X"d8", X"92", 
    X"35", X"3c", X"72", X"6c", X"63", X"2c", X"72", X"72", 
    X"63", X"2c", X"72", X"61", X"6c", X"2c", X"72", X"61", 
    X"72", X"3e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"ff", X"02", X"00", X"00", X"00", X"3b", X"0c", X"92", 
    X"b5", X"ff", X"6c", X"9e", X"95", X"03", X"01", X"04", 
    X"01", X"c1", X"21", X"e7", X"bd", X"18", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"ff", X"ff", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"ff", X"00", X"00", X"2b", X"04", X"71", 
    X"e9", X"73", X"74", X"61", X"78", X"20", X"3c", X"62", 
    X"2c", X"64", X"3e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", 
    X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"2e", X"24", 
    X"e5", X"7e", X"23", X"66", X"6f", X"7e", X"32", X"81", 
    X"0d", X"23", X"e5", X"11", X"14", X"00", X"19", X"11", 
    X"e0", X"0c", X"cd", X"4f", X"0c", X"e1", X"e5", X"11", 
    X"28", X"00", X"19", X"11", X"08", X"0d", X"cd", X"4f", 
    X"0c", X"21", X"08", X"0d", X"36", X"01", X"e1", X"e5", 
    X"11", X"4f", X"0d", X"01", X"04", X"00", X"7e", X"12", 
    X"23", X"13", X"0b", X"78", X"b1", X"c2", X"fe", X"0a", 
    X"11", X"03", X"01", X"01", X"10", X"00", X"7e", X"12", 
    X"23", X"13", X"0b", X"78", X"b1", X"c2", X"0e", X"0b", 
    X"11", X"2c", X"00", X"19", X"eb", X"0e", X"09", X"cd", 
    X"ec", X"0d", X"cd", X"92", X"0e", X"3a", X"4f", X"0d", 
    X"fe", X"76", X"ca", X"3c", X"0b", X"e6", X"df", X"fe", 
    X"dd", X"c2", X"39", X"0b", X"3a", X"50", X"0d", X"fe", 
    X"76", X"c4", X"30", X"0d", X"cd", X"8f", X"0c", X"c4", 
    X"b3", X"0c", X"e1", X"ca", X"78", X"0b", X"11", X"3c", 
    X"00", X"19", X"cd", X"53", X"0e", X"11", X"26", X"0e", 
    X"ca", X"6f", X"0b", X"11", X"2d", X"0e", X"0e", X"09", 
    X"cd", X"ec", X"0d", X"cd", X"b7", X"0d", X"11", X"48", 
    X"0e", X"0e", X"09", X"cd", X"ec", X"0d", X"21", X"ed", 
    X"0e", X"cd", X"b7", X"0d", X"11", X"50", X"0e", X"0e", 
    X"09", X"cd", X"ec", X"0d", X"e1", X"23", X"23", X"c9", 
    X"e5", X"3e", X"01", X"32", X"ee", X"0b", X"32", X"12", 
    X"0c", X"21", X"e0", X"0c", X"22", X"ef", X"0b", X"21", 
    X"08", X"0d", X"22", X"13", X"0c", X"06", X"04", X"e1", 
    X"e5", X"11", X"4f", X"0d", X"cd", X"a2", X"0b", X"06", 
    X"10", X"11", X"03", X"01", X"cd", X"a2", X"0b", X"c3", 
    X"25", X"0b", X"cd", X"ab", X"0b", X"23", X"05", X"c2", 
    X"a2", X"0b", X"c9", X"c5", X"d5", X"e5", X"4e", X"11", 
    X"14", X"00", X"19", X"7e", X"fe", X"00", X"ca", X"cc", 
    X"0b", X"06", X"08", X"0f", X"f5", X"3e", X"00", X"dc", 
    X"f1", X"0b", X"a9", X"0f", X"4f", X"f1", X"05", X"c2", 
    X"bb", X"0b", X"06", X"08", X"11", X"14", X"00", X"19", 
    X"7e", X"fe", X"00", X"ca", X"e7", X"0b", X"06", X"08", 
    X"0f", X"f5", X"3e", X"00", X"dc", X"15", X"0c", X"a9", 
    X"0f", X"4f", X"f1", X"05", X"c2", X"d8", X"0b", X"e1", 
    X"d1", X"79", X"12", X"13", X"c1", X"c9", X"00", X"00", 
    X"00", X"c5", X"e5", X"2a", X"ef", X"0b", X"46", X"21", 
    X"ee", X"0b", X"7e", X"4f", X"07", X"77", X"fe", X"01", 
    X"c2", X"0a", X"0c", X"2a", X"ef", X"0b", X"23", X"22", 
    X"ef", X"0b", X"78", X"a1", X"e1", X"c1", X"c8", X"3e", 
    X"01", X"c9", X"00", X"00", X"00", X"c5", X"e5", X"2a", 
    X"13", X"0c", X"46", X"21", X"12", X"0c", X"7e", X"4f", 
    X"07", X"77", X"fe", X"01", X"c2", X"2e", X"0c", X"2a", 
    X"13", X"0c", X"23", X"22", X"13", X"0c", X"78", X"a1", 
    X"e1", X"c1", X"c8", X"3e", X"01", X"c9", X"f5", X"c5", 
    X"d5", X"e5", X"36", X"00", X"54", X"5d", X"13", X"0b", 
    X"7e", X"12", X"23", X"13", X"0b", X"78", X"b1", X"c2", 
    X"40", X"0c", X"e1", X"d1", X"c1", X"f1", X"c9", X"d5", 
    X"eb", X"01", X"28", X"00", X"cd", X"36", X"0c", X"eb", 
    X"06", X"14", X"0e", X"01", X"16", X"00", X"5e", X"7b", 
    X"a1", X"ca", X"65", X"0c", X"14", X"79", X"07", X"4f", 
    X"fe", X"01", X"c2", X"5f", X"0c", X"23", X"05", X"c2", 
    X"5e", X"0c", X"7a", X"e6", X"f8", X"0f", X"0f", X"0f", 
    X"6f", X"26", X"00", X"7a", X"e6", X"07", X"3c", X"47", 
    X"3e", X"80", X"07", X"05", X"c2", X"82", X"0c", X"d1", 
    X"19", X"11", X"14", X"00", X"19", X"77", X"c9", X"c5", 
    X"d5", X"e5", X"21", X"e0", X"0c", X"11", X"14", X"00", 
    X"eb", X"19", X"eb", X"34", X"7e", X"fe", X"00", X"ca", 
    X"ae", X"0c", X"47", X"1a", X"a0", X"ca", X"aa", X"0c", 
    X"36", X"00", X"c1", X"d1", X"e1", X"c9", X"23", X"13", 
    X"c3", X"9b", X"0c", X"c5", X"d5", X"e5", X"21", X"08", 
    X"0d", X"11", X"14", X"00", X"eb", X"19", X"eb", X"7e", 
    X"b7", X"ca", X"db", X"0c", X"47", X"1a", X"a0", X"c2", 
    X"d7", X"0c", X"78", X"07", X"fe", X"01", X"c2", X"d5", 
    X"0c", X"36", X"00", X"23", X"13", X"77", X"af", X"e1", 
    X"d1", X"c1", X"c9", X"23", X"13", X"c3", X"bf", X"0c", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"f5", X"c5", X"d5", X"e5", X"f3", X"21", X"00", X"00", 
    X"39", X"22", X"ab", X"0d", X"31", X"05", X"01", X"e1", 
    X"e1", X"e1", X"d1", X"c1", X"f1", X"22", X"99", X"0d", 
    X"2a", X"11", X"01", X"f9", X"2a", X"99", X"0d", X"00", 
    X"00", X"00", X"00", X"22", X"99", X"0d", X"21", X"00", 
    X"00", X"da", X"60", X"0d", X"39", X"c3", X"62", X"0d", 
    X"39", X"37", X"22", X"a9", X"0d", X"2a", X"99", X"0d", 
    X"31", X"a9", X"0d", X"f5", X"c5", X"d5", X"e5", X"e5", 
    X"e5", X"2a", X"ab", X"0d", X"f9", X"fb", X"2a", X"03", 
    X"01", X"22", X"9b", X"0d", X"21", X"a7", X"0d", X"7e", 
    X"e6", X"ff", X"77", X"06", X"10", X"11", X"9b", X"0d", 
    X"21", X"ed", X"0e", X"1a", X"13", X"cd", X"6a", X"0e", 
    X"05", X"c2", X"8b", X"0d", X"e1", X"d1", X"c1", X"f1", 
    X"c9", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"7e", X"cd", X"c9", 
    X"0d", X"23", X"05", X"c2", X"ad", X"0d", X"c9", X"f5", 
    X"c5", X"e5", X"06", X"04", X"7e", X"cd", X"c9", X"0d", 
    X"23", X"05", X"c2", X"bc", X"0d", X"e1", X"c1", X"f1", 
    X"c9", X"f5", X"0f", X"0f", X"0f", X"0f", X"cd", X"d2", 
    X"0d", X"f1", X"f5", X"c5", X"d5", X"e5", X"e6", X"0f", 
    X"fe", X"0a", X"da", X"df", X"0d", X"c6", X"27", X"c6", 
    X"30", X"5f", X"0e", X"02", X"cd", X"ec", X"0d", X"e1", 
    X"d1", X"c1", X"f1", X"c9", X"f5", X"c5", X"d5", X"e5", 
    X"cd", X"05", X"00", X"e1", X"d1", X"c1", X"f1", X"c9", 
    X"38", X"30", X"38", X"30", X"20", X"69", X"6e", X"73", 
    X"74", X"72", X"75", X"63", X"74", X"69", X"6f", X"6e", 
    X"20", X"65", X"78", X"65", X"72", X"63", X"69", X"73", 
    X"65", X"72", X"0a", X"0d", X"24", X"54", X"65", X"73", 
    X"74", X"73", X"20", X"63", X"6f", X"6d", X"70", X"6c", 
    X"65", X"74", X"65", X"0a", X"0d", X"24", X"20", X"20", 
    X"4f", X"4b", X"0a", X"0d", X"24", X"20", X"20", X"45", 
    X"52", X"52", X"4f", X"52", X"20", X"2a", X"2a", X"2a", 
    X"2a", X"20", X"63", X"72", X"63", X"20", X"65", X"78", 
    X"70", X"65", X"63", X"74", X"65", X"64", X"3a", X"24", 
    X"20", X"66", X"6f", X"75", X"6e", X"64", X"3a", X"24", 
    X"0a", X"0d", X"24", X"c5", X"d5", X"e5", X"11", X"ed", 
    X"0e", X"06", X"04", X"1a", X"be", X"c2", X"66", X"0e", 
    X"23", X"13", X"05", X"c2", X"5b", X"0e", X"e1", X"d1", 
    X"c1", X"c9", X"f5", X"c5", X"d5", X"e5", X"e5", X"11", 
    X"03", X"00", X"19", X"ae", X"6f", X"26", X"00", X"29", 
    X"29", X"eb", X"21", X"f1", X"0e", X"19", X"eb", X"e1", 
    X"01", X"04", X"00", X"1a", X"a8", X"46", X"77", X"13", 
    X"23", X"0d", X"c2", X"83", X"0e", X"e1", X"d1", X"c1", 
    X"f1", X"c9", X"f5", X"c5", X"e5", X"21", X"ed", X"0e", 
    X"3e", X"ff", X"06", X"04", X"77", X"23", X"05", X"c2", 
    X"9c", X"0e", X"e1", X"c1", X"f1", X"c9", X"47", X"79", 
    X"fe", X"09", X"ca", X"d6", X"0e", X"fe", X"02", X"ca", 
    X"d2", X"0e", X"11", X"ba", X"0e", X"cd", X"d6", X"0e", 
    X"f3", X"76", X"49", X"6e", X"76", X"61", X"6c", X"69", 
    X"64", X"20", X"42", X"44", X"4f", X"53", X"20", X"66", 
    X"75", X"6e", X"63", X"74", X"69", X"6f", X"6e", X"0d", 
    X"0a", X"24", X"48", X"c3", X"e2", X"0e", X"1a", X"13", 
    X"fe", X"24", X"c8", X"4f", X"cd", X"e2", X"0e", X"c3", 
    X"d6", X"0e", X"db", X"81", X"e6", X"01", X"ca", X"e2", 
    X"0e", X"79", X"d3", X"80", X"c9", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"77", X"07", X"30", 
    X"96", X"ee", X"0e", X"61", X"2c", X"99", X"09", X"51", 
    X"ba", X"07", X"6d", X"c4", X"19", X"70", X"6a", X"f4", 
    X"8f", X"e9", X"63", X"a5", X"35", X"9e", X"64", X"95", 
    X"a3", X"0e", X"db", X"88", X"32", X"79", X"dc", X"b8", 
    X"a4", X"e0", X"d5", X"e9", X"1e", X"97", X"d2", X"d9", 
    X"88", X"09", X"b6", X"4c", X"2b", X"7e", X"b1", X"7c", 
    X"bd", X"e7", X"b8", X"2d", X"07", X"90", X"bf", X"1d", 
    X"91", X"1d", X"b7", X"10", X"64", X"6a", X"b0", X"20", 
    X"f2", X"f3", X"b9", X"71", X"48", X"84", X"be", X"41", 
    X"de", X"1a", X"da", X"d4", X"7d", X"6d", X"dd", X"e4", 
    X"eb", X"f4", X"d4", X"b5", X"51", X"83", X"d3", X"85", 
    X"c7", X"13", X"6c", X"98", X"56", X"64", X"6b", X"a8", 
    X"c0", X"fd", X"62", X"f9", X"7a", X"8a", X"65", X"c9", 
    X"ec", X"14", X"01", X"5c", X"4f", X"63", X"06", X"6c", 
    X"d9", X"fa", X"0f", X"3d", X"63", X"8d", X"08", X"0d", 
    X"f5", X"3b", X"6e", X"20", X"c8", X"4c", X"69", X"10", 
    X"5e", X"d5", X"60", X"41", X"e4", X"a2", X"67", X"71", 
    X"72", X"3c", X"03", X"e4", X"d1", X"4b", X"04", X"d4", 
    X"47", X"d2", X"0d", X"85", X"fd", X"a5", X"0a", X"b5", 
    X"6b", X"35", X"b5", X"a8", X"fa", X"42", X"b2", X"98", 
    X"6c", X"db", X"bb", X"c9", X"d6", X"ac", X"bc", X"f9", 
    X"40", X"32", X"d8", X"6c", X"e3", X"45", X"df", X"5c", 
    X"75", X"dc", X"d6", X"0d", X"cf", X"ab", X"d1", X"3d", 
    X"59", X"26", X"d9", X"30", X"ac", X"51", X"de", X"00", 
    X"3a", X"c8", X"d7", X"51", X"80", X"bf", X"d0", X"61", 
    X"16", X"21", X"b4", X"f4", X"b5", X"56", X"b3", X"c4", 
    X"23", X"cf", X"ba", X"95", X"99", X"b8", X"bd", X"a5", 
    X"0f", X"28", X"02", X"b8", X"9e", X"5f", X"05", X"88", 
    X"08", X"c6", X"0c", X"d9", X"b2", X"b1", X"0b", X"e9", 
    X"24", X"2f", X"6f", X"7c", X"87", X"58", X"68", X"4c", 
    X"11", X"c1", X"61", X"1d", X"ab", X"b6", X"66", X"2d", 
    X"3d", X"76", X"dc", X"41", X"90", X"01", X"db", X"71", 
    X"06", X"98", X"d2", X"20", X"bc", X"ef", X"d5", X"10", 
    X"2a", X"71", X"b1", X"85", X"89", X"06", X"b6", X"b5", 
    X"1f", X"9f", X"bf", X"e4", X"a5", X"e8", X"b8", X"d4", 
    X"33", X"78", X"07", X"c9", X"a2", X"0f", X"00", X"f9", 
    X"34", X"96", X"09", X"a8", X"8e", X"e1", X"0e", X"98", 
    X"18", X"7f", X"6a", X"0d", X"bb", X"08", X"6d", X"3d", 
    X"2d", X"91", X"64", X"6c", X"97", X"e6", X"63", X"5c", 
    X"01", X"6b", X"6b", X"51", X"f4", X"1c", X"6c", X"61", 
    X"62", X"85", X"65", X"30", X"d8", X"f2", X"62", X"00", 
    X"4e", X"6c", X"06", X"95", X"ed", X"1b", X"01", X"a5", 
    X"7b", X"82", X"08", X"f4", X"c1", X"f5", X"0f", X"c4", 
    X"57", X"65", X"b0", X"d9", X"c6", X"12", X"b7", X"e9", 
    X"50", X"8b", X"be", X"b8", X"ea", X"fc", X"b9", X"88", 
    X"7c", X"62", X"dd", X"1d", X"df", X"15", X"da", X"2d", 
    X"49", X"8c", X"d3", X"7c", X"f3", X"fb", X"d4", X"4c", 
    X"65", X"4d", X"b2", X"61", X"58", X"3a", X"b5", X"51", 
    X"ce", X"a3", X"bc", X"00", X"74", X"d4", X"bb", X"30", 
    X"e2", X"4a", X"df", X"a5", X"41", X"3d", X"d8", X"95", 
    X"d7", X"a4", X"d1", X"c4", X"6d", X"d3", X"d6", X"f4", 
    X"fb", X"43", X"69", X"e9", X"6a", X"34", X"6e", X"d9", 
    X"fc", X"ad", X"67", X"88", X"46", X"da", X"60", X"b8", 
    X"d0", X"44", X"04", X"2d", X"73", X"33", X"03", X"1d", 
    X"e5", X"aa", X"0a", X"4c", X"5f", X"dd", X"0d", X"7c", 
    X"c9", X"50", X"05", X"71", X"3c", X"27", X"02", X"41", 
    X"aa", X"be", X"0b", X"10", X"10", X"c9", X"0c", X"20", 
    X"86", X"57", X"68", X"b5", X"25", X"20", X"6f", X"85", 
    X"b3", X"b9", X"66", X"d4", X"09", X"ce", X"61", X"e4", 
    X"9f", X"5e", X"de", X"f9", X"0e", X"29", X"d9", X"c9", 
    X"98", X"b0", X"d0", X"98", X"22", X"c7", X"d7", X"a8", 
    X"b4", X"59", X"b3", X"3d", X"17", X"2e", X"b4", X"0d", 
    X"81", X"b7", X"bd", X"5c", X"3b", X"c0", X"ba", X"6c", 
    X"ad", X"ed", X"b8", X"83", X"20", X"9a", X"bf", X"b3", 
    X"b6", X"03", X"b6", X"e2", X"0c", X"74", X"b1", X"d2", 
    X"9a", X"ea", X"d5", X"47", X"39", X"9d", X"d2", X"77", 
    X"af", X"04", X"db", X"26", X"15", X"73", X"dc", X"16", 
    X"83", X"e3", X"63", X"0b", X"12", X"94", X"64", X"3b", 
    X"84", X"0d", X"6d", X"6a", X"3e", X"7a", X"6a", X"5a", 
    X"a8", X"e4", X"0e", X"cf", X"0b", X"93", X"09", X"ff", 
    X"9d", X"0a", X"00", X"ae", X"27", X"7d", X"07", X"9e", 
    X"b1", X"f0", X"0f", X"93", X"44", X"87", X"08", X"a3", 
    X"d2", X"1e", X"01", X"f2", X"68", X"69", X"06", X"c2", 
    X"fe", X"f7", X"62", X"57", X"5d", X"80", X"65", X"67", 
    X"cb", X"19", X"6c", X"36", X"71", X"6e", X"6b", X"06", 
    X"e7", X"fe", X"d4", X"1b", X"76", X"89", X"d3", X"2b", 
    X"e0", X"10", X"da", X"7a", X"5a", X"67", X"dd", X"4a", 
    X"cc", X"f9", X"b9", X"df", X"6f", X"8e", X"be", X"ef", 
    X"f9", X"17", X"b7", X"be", X"43", X"60", X"b0", X"8e", 
    X"d5", X"d6", X"d6", X"a3", X"e8", X"a1", X"d1", X"93", 
    X"7e", X"38", X"d8", X"c2", X"c4", X"4f", X"df", X"f2", 
    X"52", X"d1", X"bb", X"67", X"f1", X"a6", X"bc", X"57", 
    X"67", X"3f", X"b5", X"06", X"dd", X"48", X"b2", X"36", 
    X"4b", X"d8", X"0d", X"2b", X"da", X"af", X"0a", X"1b", 
    X"4c", X"36", X"03", X"4a", X"f6", X"41", X"04", X"7a", 
    X"60", X"df", X"60", X"ef", X"c3", X"a8", X"67", X"df", 
    X"55", X"31", X"6e", X"8e", X"ef", X"46", X"69", X"be", 
    X"79", X"cb", X"61", X"b3", X"8c", X"bc", X"66", X"83", 
    X"1a", X"25", X"6f", X"d2", X"a0", X"52", X"68", X"e2", 
    X"36", X"cc", X"0c", X"77", X"95", X"bb", X"0b", X"47", 
    X"03", X"22", X"02", X"16", X"b9", X"55", X"05", X"26", 
    X"2f", X"c5", X"ba", X"3b", X"be", X"b2", X"bd", X"0b", 
    X"28", X"2b", X"b4", X"5a", X"92", X"5c", X"b3", X"6a", 
    X"04", X"c2", X"d7", X"ff", X"a7", X"b5", X"d0", X"cf", 
    X"31", X"2c", X"d9", X"9e", X"8b", X"5b", X"de", X"ae", 
    X"1d", X"9b", X"64", X"c2", X"b0", X"ec", X"63", X"f2", 
    X"26", X"75", X"6a", X"a3", X"9c", X"02", X"6d", X"93", 
    X"0a", X"9c", X"09", X"06", X"a9", X"eb", X"0e", X"36", 
    X"3f", X"72", X"07", X"67", X"85", X"05", X"00", X"57", 
    X"13", X"95", X"bf", X"4a", X"82", X"e2", X"b8", X"7a", 
    X"14", X"7b", X"b1", X"2b", X"ae", X"0c", X"b6", X"1b", 
    X"38", X"92", X"d2", X"8e", X"9b", X"e5", X"d5", X"be", 
    X"0d", X"7c", X"dc", X"ef", X"b7", X"0b", X"db", X"df", 
    X"21", X"86", X"d3", X"d2", X"d4", X"f1", X"d4", X"e2", 
    X"42", X"68", X"dd", X"b3", X"f8", X"1f", X"da", X"83", 
    X"6e", X"81", X"be", X"16", X"cd", X"f6", X"b9", X"26", 
    X"5b", X"6f", X"b0", X"77", X"e1", X"18", X"b7", X"47", 
    X"77", X"88", X"08", X"5a", X"e6", X"ff", X"0f", X"6a", 
    X"70", X"66", X"06", X"3b", X"ca", X"11", X"01", X"0b", 
    X"5c", X"8f", X"65", X"9e", X"ff", X"f8", X"62", X"ae", 
    X"69", X"61", X"6b", X"ff", X"d3", X"16", X"6c", X"cf", 
    X"45", X"a0", X"0a", X"e2", X"78", X"d7", X"0d", X"d2", 
    X"ee", X"4e", X"04", X"83", X"54", X"39", X"03", X"b3", 
    X"c2", X"a7", X"67", X"26", X"61", X"d0", X"60", X"16", 
    X"f7", X"49", X"69", X"47", X"4d", X"3e", X"6e", X"77", 
    X"db", X"ae", X"d1", X"6a", X"4a", X"d9", X"d6", X"5a", 
    X"dc", X"40", X"df", X"0b", X"66", X"37", X"d8", X"3b", 
    X"f0", X"a9", X"bc", X"ae", X"53", X"de", X"bb", X"9e", 
    X"c5", X"47", X"b2", X"cf", X"7f", X"30", X"b5", X"ff", 
    X"e9", X"bd", X"bd", X"f2", X"1c", X"ca", X"ba", X"c2", 
    X"8a", X"53", X"b3", X"93", X"30", X"24", X"b4", X"a3", 
    X"a6", X"ba", X"d0", X"36", X"05", X"cd", X"d7", X"06", 
    X"93", X"54", X"de", X"57", X"29", X"23", X"d9", X"67", 
    X"bf", X"b3", X"66", X"7a", X"2e", X"c4", X"61", X"4a", 
    X"b8", X"5d", X"68", X"1b", X"02", X"2a", X"6f", X"2b", 
    X"94", X"b4", X"0b", X"be", X"37", X"c3", X"0c", X"8e", 
    X"a1", X"5a", X"05", X"df", X"1b", X"2d", X"02", X"ef", 
    X"8d" 
);

end package obj_code_pkg;
