-----------------------------------------------------------------
--                                                             --
-----------------------------------------------------------------
--                                                             --
-- Copyright (C) 2013 Stefano Tonello                          --
--                                                             --
-- This source file may be used and distributed without        --
-- restriction provided that this copyright statement is not   --
-- removed from the file and that any derivative work contains --
-- the original copyright notice and the associated disclaimer.--
--                                                             --
-- THIS SOFTWARE IS PROVIDED ``AS IS'' AND WITHOUT ANY         --
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   --
-- TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS   --
-- FOR A PARTICULAR PURPOSE. IN NO EVENT SHALL THE AUTHOR      --
-- OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,         --
-- INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES    --
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE   --
-- GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR        --
-- BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF  --
-- LIABILITY, WHETHER IN  CONTRACT, STRICT LIABILITY, OR TORT  --
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT  --
-- OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE         --
-- POSSIBILITY OF SUCH DAMAGE.                                 --
--                                                             --
-----------------------------------------------------------------

---------------------------------------------------------------
-- G.729a ASIP Constant Data ROM content
---------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library WORK;
use work.G729A_ASIP_PKG.all;
use work.G729A_ASIP_CFG_PKG.all;

package G729A_ASIP_ROMD_PKG is

--WIDTH=16;
--DEPTH=3072;

--ADDRESS_RADIX=UNS;
--DATA_RADIX=DEC;

--CONTENT BEGIN

  subtype ROMD_WORD_T is std_logic_vector(SDLEN-1 downto 0);

  type ROMD_DATA_T is array (0 to CMEM_LIMIT-1) of ROMD_WORD_T;

  constant ROMD_INIT_DATA : ROMD_DATA_T := (

    to_std_logic_vector(to_signed(2621,SDLEN)),
    to_std_logic_vector(to_signed(2623,SDLEN)),
    to_std_logic_vector(to_signed(2629,SDLEN)),
    to_std_logic_vector(to_signed(2638,SDLEN)),
    to_std_logic_vector(to_signed(2651,SDLEN)),
    to_std_logic_vector(to_signed(2668,SDLEN)),
    to_std_logic_vector(to_signed(2689,SDLEN)),
    to_std_logic_vector(to_signed(2713,SDLEN)),
    to_std_logic_vector(to_signed(2741,SDLEN)),
    to_std_logic_vector(to_signed(2772,SDLEN)),
    to_std_logic_vector(to_signed(2808,SDLEN)),
    to_std_logic_vector(to_signed(2847,SDLEN)),
    to_std_logic_vector(to_signed(2890,SDLEN)),
    to_std_logic_vector(to_signed(2936,SDLEN)),
    to_std_logic_vector(to_signed(2986,SDLEN)),
    to_std_logic_vector(to_signed(3040,SDLEN)),
    to_std_logic_vector(to_signed(3097,SDLEN)),
    to_std_logic_vector(to_signed(3158,SDLEN)),
    to_std_logic_vector(to_signed(3223,SDLEN)),
    to_std_logic_vector(to_signed(3291,SDLEN)),
    to_std_logic_vector(to_signed(3363,SDLEN)),
    to_std_logic_vector(to_signed(3438,SDLEN)),
    to_std_logic_vector(to_signed(3517,SDLEN)),
    to_std_logic_vector(to_signed(3599,SDLEN)),
    to_std_logic_vector(to_signed(3685,SDLEN)),
    to_std_logic_vector(to_signed(3774,SDLEN)),
    to_std_logic_vector(to_signed(3867,SDLEN)),
    to_std_logic_vector(to_signed(3963,SDLEN)),
    to_std_logic_vector(to_signed(4063,SDLEN)),
    to_std_logic_vector(to_signed(4166,SDLEN)),
    to_std_logic_vector(to_signed(4272,SDLEN)),
    to_std_logic_vector(to_signed(4382,SDLEN)),
    to_std_logic_vector(to_signed(4495,SDLEN)),
    to_std_logic_vector(to_signed(4611,SDLEN)),
    to_std_logic_vector(to_signed(4731,SDLEN)),
    to_std_logic_vector(to_signed(4853,SDLEN)),
    to_std_logic_vector(to_signed(4979,SDLEN)),
    to_std_logic_vector(to_signed(5108,SDLEN)),
    to_std_logic_vector(to_signed(5240,SDLEN)),
    to_std_logic_vector(to_signed(5376,SDLEN)),
    to_std_logic_vector(to_signed(5514,SDLEN)),
    to_std_logic_vector(to_signed(5655,SDLEN)),
    to_std_logic_vector(to_signed(5800,SDLEN)),
    to_std_logic_vector(to_signed(5947,SDLEN)),
    to_std_logic_vector(to_signed(6097,SDLEN)),
    to_std_logic_vector(to_signed(6250,SDLEN)),
    to_std_logic_vector(to_signed(6406,SDLEN)),
    to_std_logic_vector(to_signed(6565,SDLEN)),
    to_std_logic_vector(to_signed(6726,SDLEN)),
    to_std_logic_vector(to_signed(6890,SDLEN)),
    to_std_logic_vector(to_signed(7057,SDLEN)),
    to_std_logic_vector(to_signed(7227,SDLEN)),
    to_std_logic_vector(to_signed(7399,SDLEN)),
    to_std_logic_vector(to_signed(7573,SDLEN)),
    to_std_logic_vector(to_signed(7750,SDLEN)),
    to_std_logic_vector(to_signed(7930,SDLEN)),
    to_std_logic_vector(to_signed(8112,SDLEN)),
    to_std_logic_vector(to_signed(8296,SDLEN)),
    to_std_logic_vector(to_signed(8483,SDLEN)),
    to_std_logic_vector(to_signed(8672,SDLEN)),
    to_std_logic_vector(to_signed(8863,SDLEN)),
    to_std_logic_vector(to_signed(9057,SDLEN)),
    to_std_logic_vector(to_signed(9252,SDLEN)),
    to_std_logic_vector(to_signed(9450,SDLEN)),
    to_std_logic_vector(to_signed(9650,SDLEN)),
    to_std_logic_vector(to_signed(9852,SDLEN)),
    to_std_logic_vector(to_signed(10055,SDLEN)),
    to_std_logic_vector(to_signed(10261,SDLEN)),
    to_std_logic_vector(to_signed(10468,SDLEN)),
    to_std_logic_vector(to_signed(10677,SDLEN)),
    to_std_logic_vector(to_signed(10888,SDLEN)),
    to_std_logic_vector(to_signed(11101,SDLEN)),
    to_std_logic_vector(to_signed(11315,SDLEN)),
    to_std_logic_vector(to_signed(11531,SDLEN)),
    to_std_logic_vector(to_signed(11748,SDLEN)),
    to_std_logic_vector(to_signed(11967,SDLEN)),
    to_std_logic_vector(to_signed(12187,SDLEN)),
    to_std_logic_vector(to_signed(12409,SDLEN)),
    to_std_logic_vector(to_signed(12632,SDLEN)),
    to_std_logic_vector(to_signed(12856,SDLEN)),
    to_std_logic_vector(to_signed(13082,SDLEN)),
    to_std_logic_vector(to_signed(13308,SDLEN)),
    to_std_logic_vector(to_signed(13536,SDLEN)),
    to_std_logic_vector(to_signed(13764,SDLEN)),
    to_std_logic_vector(to_signed(13994,SDLEN)),
    to_std_logic_vector(to_signed(14225,SDLEN)),
    to_std_logic_vector(to_signed(14456,SDLEN)),
    to_std_logic_vector(to_signed(14688,SDLEN)),
    to_std_logic_vector(to_signed(14921,SDLEN)),
    to_std_logic_vector(to_signed(15155,SDLEN)),
    to_std_logic_vector(to_signed(15389,SDLEN)),
    to_std_logic_vector(to_signed(15624,SDLEN)),
    to_std_logic_vector(to_signed(15859,SDLEN)),
    to_std_logic_vector(to_signed(16095,SDLEN)),
    to_std_logic_vector(to_signed(16331,SDLEN)),
    to_std_logic_vector(to_signed(16568,SDLEN)),
    to_std_logic_vector(to_signed(16805,SDLEN)),
    to_std_logic_vector(to_signed(17042,SDLEN)),
    to_std_logic_vector(to_signed(17279,SDLEN)),
    to_std_logic_vector(to_signed(17516,SDLEN)),
    to_std_logic_vector(to_signed(17754,SDLEN)),
    to_std_logic_vector(to_signed(17991,SDLEN)),
    to_std_logic_vector(to_signed(18228,SDLEN)),
    to_std_logic_vector(to_signed(18465,SDLEN)),
    to_std_logic_vector(to_signed(18702,SDLEN)),
    to_std_logic_vector(to_signed(18939,SDLEN)),
    to_std_logic_vector(to_signed(19175,SDLEN)),
    to_std_logic_vector(to_signed(19411,SDLEN)),
    to_std_logic_vector(to_signed(19647,SDLEN)),
    to_std_logic_vector(to_signed(19882,SDLEN)),
    to_std_logic_vector(to_signed(20117,SDLEN)),
    to_std_logic_vector(to_signed(20350,SDLEN)),
    to_std_logic_vector(to_signed(20584,SDLEN)),
    to_std_logic_vector(to_signed(20816,SDLEN)),
    to_std_logic_vector(to_signed(21048,SDLEN)),
    to_std_logic_vector(to_signed(21279,SDLEN)),
    to_std_logic_vector(to_signed(21509,SDLEN)),
    to_std_logic_vector(to_signed(21738,SDLEN)),
    to_std_logic_vector(to_signed(21967,SDLEN)),
    to_std_logic_vector(to_signed(22194,SDLEN)),
    to_std_logic_vector(to_signed(22420,SDLEN)),
    to_std_logic_vector(to_signed(22644,SDLEN)),
    to_std_logic_vector(to_signed(22868,SDLEN)),
    to_std_logic_vector(to_signed(23090,SDLEN)),
    to_std_logic_vector(to_signed(23311,SDLEN)),
    to_std_logic_vector(to_signed(23531,SDLEN)),
    to_std_logic_vector(to_signed(23749,SDLEN)),
    to_std_logic_vector(to_signed(23965,SDLEN)),
    to_std_logic_vector(to_signed(24181,SDLEN)),
    to_std_logic_vector(to_signed(24394,SDLEN)),
    to_std_logic_vector(to_signed(24606,SDLEN)),
    to_std_logic_vector(to_signed(24816,SDLEN)),
    to_std_logic_vector(to_signed(25024,SDLEN)),
    to_std_logic_vector(to_signed(25231,SDLEN)),
    to_std_logic_vector(to_signed(25435,SDLEN)),
    to_std_logic_vector(to_signed(25638,SDLEN)),
    to_std_logic_vector(to_signed(25839,SDLEN)),
    to_std_logic_vector(to_signed(26037,SDLEN)),
    to_std_logic_vector(to_signed(26234,SDLEN)),
    to_std_logic_vector(to_signed(26428,SDLEN)),
    to_std_logic_vector(to_signed(26621,SDLEN)),
    to_std_logic_vector(to_signed(26811,SDLEN)),
    to_std_logic_vector(to_signed(26999,SDLEN)),
    to_std_logic_vector(to_signed(27184,SDLEN)),
    to_std_logic_vector(to_signed(27368,SDLEN)),
    to_std_logic_vector(to_signed(27548,SDLEN)),
    to_std_logic_vector(to_signed(27727,SDLEN)),
    to_std_logic_vector(to_signed(27903,SDLEN)),
    to_std_logic_vector(to_signed(28076,SDLEN)),
    to_std_logic_vector(to_signed(28247,SDLEN)),
    to_std_logic_vector(to_signed(28415,SDLEN)),
    to_std_logic_vector(to_signed(28581,SDLEN)),
    to_std_logic_vector(to_signed(28743,SDLEN)),
    to_std_logic_vector(to_signed(28903,SDLEN)),
    to_std_logic_vector(to_signed(29061,SDLEN)),
    to_std_logic_vector(to_signed(29215,SDLEN)),
    to_std_logic_vector(to_signed(29367,SDLEN)),
    to_std_logic_vector(to_signed(29515,SDLEN)),
    to_std_logic_vector(to_signed(29661,SDLEN)),
    to_std_logic_vector(to_signed(29804,SDLEN)),
    to_std_logic_vector(to_signed(29944,SDLEN)),
    to_std_logic_vector(to_signed(30081,SDLEN)),
    to_std_logic_vector(to_signed(30214,SDLEN)),
    to_std_logic_vector(to_signed(30345,SDLEN)),
    to_std_logic_vector(to_signed(30472,SDLEN)),
    to_std_logic_vector(to_signed(30597,SDLEN)),
    to_std_logic_vector(to_signed(30718,SDLEN)),
    to_std_logic_vector(to_signed(30836,SDLEN)),
    to_std_logic_vector(to_signed(30950,SDLEN)),
    to_std_logic_vector(to_signed(31062,SDLEN)),
    to_std_logic_vector(to_signed(31170,SDLEN)),
    to_std_logic_vector(to_signed(31274,SDLEN)),
    to_std_logic_vector(to_signed(31376,SDLEN)),
    to_std_logic_vector(to_signed(31474,SDLEN)),
    to_std_logic_vector(to_signed(31568,SDLEN)),
    to_std_logic_vector(to_signed(31659,SDLEN)),
    to_std_logic_vector(to_signed(31747,SDLEN)),
    to_std_logic_vector(to_signed(31831,SDLEN)),
    to_std_logic_vector(to_signed(31911,SDLEN)),
    to_std_logic_vector(to_signed(31988,SDLEN)),
    to_std_logic_vector(to_signed(32062,SDLEN)),
    to_std_logic_vector(to_signed(32132,SDLEN)),
    to_std_logic_vector(to_signed(32198,SDLEN)),
    to_std_logic_vector(to_signed(32261,SDLEN)),
    to_std_logic_vector(to_signed(32320,SDLEN)),
    to_std_logic_vector(to_signed(32376,SDLEN)),
    to_std_logic_vector(to_signed(32428,SDLEN)),
    to_std_logic_vector(to_signed(32476,SDLEN)),
    to_std_logic_vector(to_signed(32521,SDLEN)),
    to_std_logic_vector(to_signed(32561,SDLEN)),
    to_std_logic_vector(to_signed(32599,SDLEN)),
    to_std_logic_vector(to_signed(32632,SDLEN)),
    to_std_logic_vector(to_signed(32662,SDLEN)),
    to_std_logic_vector(to_signed(32688,SDLEN)),
    to_std_logic_vector(to_signed(32711,SDLEN)),
    to_std_logic_vector(to_signed(32729,SDLEN)),
    to_std_logic_vector(to_signed(32744,SDLEN)),
    to_std_logic_vector(to_signed(32755,SDLEN)),
    to_std_logic_vector(to_signed(32763,SDLEN)),
    to_std_logic_vector(to_signed(32767,SDLEN)),
    to_std_logic_vector(to_signed(32767,SDLEN)),
    to_std_logic_vector(to_signed(32741,SDLEN)),
    to_std_logic_vector(to_signed(32665,SDLEN)),
    to_std_logic_vector(to_signed(32537,SDLEN)),
    to_std_logic_vector(to_signed(32359,SDLEN)),
    to_std_logic_vector(to_signed(32129,SDLEN)),
    to_std_logic_vector(to_signed(31850,SDLEN)),
    to_std_logic_vector(to_signed(31521,SDLEN)),
    to_std_logic_vector(to_signed(31143,SDLEN)),
    to_std_logic_vector(to_signed(30716,SDLEN)),
    to_std_logic_vector(to_signed(30242,SDLEN)),
    to_std_logic_vector(to_signed(29720,SDLEN)),
    to_std_logic_vector(to_signed(29151,SDLEN)),
    to_std_logic_vector(to_signed(28538,SDLEN)),
    to_std_logic_vector(to_signed(27879,SDLEN)),
    to_std_logic_vector(to_signed(27177,SDLEN)),
    to_std_logic_vector(to_signed(26433,SDLEN)),
    to_std_logic_vector(to_signed(25647,SDLEN)),
    to_std_logic_vector(to_signed(24821,SDLEN)),
    to_std_logic_vector(to_signed(23957,SDLEN)),
    to_std_logic_vector(to_signed(23055,SDLEN)),
    to_std_logic_vector(to_signed(22117,SDLEN)),
    to_std_logic_vector(to_signed(21145,SDLEN)),
    to_std_logic_vector(to_signed(20139,SDLEN)),
    to_std_logic_vector(to_signed(19102,SDLEN)),
    to_std_logic_vector(to_signed(18036,SDLEN)),
    to_std_logic_vector(to_signed(16941,SDLEN)),
    to_std_logic_vector(to_signed(15820,SDLEN)),
    to_std_logic_vector(to_signed(14674,SDLEN)),
    to_std_logic_vector(to_signed(13505,SDLEN)),
    to_std_logic_vector(to_signed(12315,SDLEN)),
    to_std_logic_vector(to_signed(11106,SDLEN)),
    to_std_logic_vector(to_signed(9879,SDLEN)),
    to_std_logic_vector(to_signed(8637,SDLEN)),
    to_std_logic_vector(to_signed(7381,SDLEN)),
    to_std_logic_vector(to_signed(6114,SDLEN)),
    to_std_logic_vector(to_signed(4838,SDLEN)),
    to_std_logic_vector(to_signed(3554,SDLEN)),
    to_std_logic_vector(to_signed(2264,SDLEN)),
    to_std_logic_vector(to_signed(971,SDLEN)),
    to_std_logic_vector(to_signed(32728,SDLEN)),
    to_std_logic_vector(to_signed(32619,SDLEN)),
    to_std_logic_vector(to_signed(32438,SDLEN)),
    to_std_logic_vector(to_signed(32187,SDLEN)),
    to_std_logic_vector(to_signed(31867,SDLEN)),
    to_std_logic_vector(to_signed(31480,SDLEN)),
    to_std_logic_vector(to_signed(31029,SDLEN)),
    to_std_logic_vector(to_signed(30517,SDLEN)),
    to_std_logic_vector(to_signed(29946,SDLEN)),
    to_std_logic_vector(to_signed(29321,SDLEN)),
    to_std_logic_vector(to_signed(11904,SDLEN)),
    to_std_logic_vector(to_signed(17280,SDLEN)),
    to_std_logic_vector(to_signed(30720,SDLEN)),
    to_std_logic_vector(to_signed(25856,SDLEN)),
    to_std_logic_vector(to_signed(24192,SDLEN)),
    to_std_logic_vector(to_signed(28992,SDLEN)),
    to_std_logic_vector(to_signed(24384,SDLEN)),
    to_std_logic_vector(to_signed(7360,SDLEN)),
    to_std_logic_vector(to_signed(19520,SDLEN)),
    to_std_logic_vector(to_signed(14784,SDLEN)),
    to_std_logic_vector(to_signed(32767,SDLEN)),
    to_std_logic_vector(to_signed(32729,SDLEN)),
    to_std_logic_vector(to_signed(32610,SDLEN)),
    to_std_logic_vector(to_signed(32413,SDLEN)),
    to_std_logic_vector(to_signed(32138,SDLEN)),
    to_std_logic_vector(to_signed(31786,SDLEN)),
    to_std_logic_vector(to_signed(31357,SDLEN)),
    to_std_logic_vector(to_signed(30853,SDLEN)),
    to_std_logic_vector(to_signed(30274,SDLEN)),
    to_std_logic_vector(to_signed(29622,SDLEN)),
    to_std_logic_vector(to_signed(28899,SDLEN)),
    to_std_logic_vector(to_signed(28106,SDLEN)),
    to_std_logic_vector(to_signed(27246,SDLEN)),
    to_std_logic_vector(to_signed(26320,SDLEN)),
    to_std_logic_vector(to_signed(25330,SDLEN)),
    to_std_logic_vector(to_signed(24279,SDLEN)),
    to_std_logic_vector(to_signed(23170,SDLEN)),
    to_std_logic_vector(to_signed(22006,SDLEN)),
    to_std_logic_vector(to_signed(20788,SDLEN)),
    to_std_logic_vector(to_signed(19520,SDLEN)),
    to_std_logic_vector(to_signed(18205,SDLEN)),
    to_std_logic_vector(to_signed(16846,SDLEN)),
    to_std_logic_vector(to_signed(15447,SDLEN)),
    to_std_logic_vector(to_signed(14010,SDLEN)),
    to_std_logic_vector(to_signed(12540,SDLEN)),
    to_std_logic_vector(to_signed(11039,SDLEN)),
    to_std_logic_vector(to_signed(9512,SDLEN)),
    to_std_logic_vector(to_signed(7962,SDLEN)),
    to_std_logic_vector(to_signed(6393,SDLEN)),
    to_std_logic_vector(to_signed(4808,SDLEN)),
    to_std_logic_vector(to_signed(3212,SDLEN)),
    to_std_logic_vector(to_signed(1608,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(-1608,SDLEN)),
    to_std_logic_vector(to_signed(-3212,SDLEN)),
    to_std_logic_vector(to_signed(-4808,SDLEN)),
    to_std_logic_vector(to_signed(-6393,SDLEN)),
    to_std_logic_vector(to_signed(-7962,SDLEN)),
    to_std_logic_vector(to_signed(-9512,SDLEN)),
    to_std_logic_vector(to_signed(-11039,SDLEN)),
    to_std_logic_vector(to_signed(-12540,SDLEN)),
    to_std_logic_vector(to_signed(-14010,SDLEN)),
    to_std_logic_vector(to_signed(-15447,SDLEN)),
    to_std_logic_vector(to_signed(-16846,SDLEN)),
    to_std_logic_vector(to_signed(-18205,SDLEN)),
    to_std_logic_vector(to_signed(-19520,SDLEN)),
    to_std_logic_vector(to_signed(-20788,SDLEN)),
    to_std_logic_vector(to_signed(-22006,SDLEN)),
    to_std_logic_vector(to_signed(-23170,SDLEN)),
    to_std_logic_vector(to_signed(-24279,SDLEN)),
    to_std_logic_vector(to_signed(-25330,SDLEN)),
    to_std_logic_vector(to_signed(-26320,SDLEN)),
    to_std_logic_vector(to_signed(-27246,SDLEN)),
    to_std_logic_vector(to_signed(-28106,SDLEN)),
    to_std_logic_vector(to_signed(-28899,SDLEN)),
    to_std_logic_vector(to_signed(-29622,SDLEN)),
    to_std_logic_vector(to_signed(-30274,SDLEN)),
    to_std_logic_vector(to_signed(-30853,SDLEN)),
    to_std_logic_vector(to_signed(-31357,SDLEN)),
    to_std_logic_vector(to_signed(-31786,SDLEN)),
    to_std_logic_vector(to_signed(-32138,SDLEN)),
    to_std_logic_vector(to_signed(-32413,SDLEN)),
    to_std_logic_vector(to_signed(-32610,SDLEN)),
    to_std_logic_vector(to_signed(-32729,SDLEN)),
    to_std_logic_vector(to_signed(-32768,SDLEN)),
    to_std_logic_vector(to_signed(-26887,SDLEN)),
    to_std_logic_vector(to_signed(-8812,SDLEN)),
    to_std_logic_vector(to_signed(-5323,SDLEN)),
    to_std_logic_vector(to_signed(-3813,SDLEN)),
    to_std_logic_vector(to_signed(-2979,SDLEN)),
    to_std_logic_vector(to_signed(-2444,SDLEN)),
    to_std_logic_vector(to_signed(-2081,SDLEN)),
    to_std_logic_vector(to_signed(-1811,SDLEN)),
    to_std_logic_vector(to_signed(-1608,SDLEN)),
    to_std_logic_vector(to_signed(-1450,SDLEN)),
    to_std_logic_vector(to_signed(-1322,SDLEN)),
    to_std_logic_vector(to_signed(-1219,SDLEN)),
    to_std_logic_vector(to_signed(-1132,SDLEN)),
    to_std_logic_vector(to_signed(-1059,SDLEN)),
    to_std_logic_vector(to_signed(-998,SDLEN)),
    to_std_logic_vector(to_signed(-946,SDLEN)),
    to_std_logic_vector(to_signed(-901,SDLEN)),
    to_std_logic_vector(to_signed(-861,SDLEN)),
    to_std_logic_vector(to_signed(-827,SDLEN)),
    to_std_logic_vector(to_signed(-797,SDLEN)),
    to_std_logic_vector(to_signed(-772,SDLEN)),
    to_std_logic_vector(to_signed(-750,SDLEN)),
    to_std_logic_vector(to_signed(-730,SDLEN)),
    to_std_logic_vector(to_signed(-713,SDLEN)),
    to_std_logic_vector(to_signed(-699,SDLEN)),
    to_std_logic_vector(to_signed(-687,SDLEN)),
    to_std_logic_vector(to_signed(-677,SDLEN)),
    to_std_logic_vector(to_signed(-668,SDLEN)),
    to_std_logic_vector(to_signed(-662,SDLEN)),
    to_std_logic_vector(to_signed(-657,SDLEN)),
    to_std_logic_vector(to_signed(-654,SDLEN)),
    to_std_logic_vector(to_signed(-652,SDLEN)),
    to_std_logic_vector(to_signed(-652,SDLEN)),
    to_std_logic_vector(to_signed(-654,SDLEN)),
    to_std_logic_vector(to_signed(-657,SDLEN)),
    to_std_logic_vector(to_signed(-662,SDLEN)),
    to_std_logic_vector(to_signed(-668,SDLEN)),
    to_std_logic_vector(to_signed(-677,SDLEN)),
    to_std_logic_vector(to_signed(-687,SDLEN)),
    to_std_logic_vector(to_signed(-699,SDLEN)),
    to_std_logic_vector(to_signed(-713,SDLEN)),
    to_std_logic_vector(to_signed(-730,SDLEN)),
    to_std_logic_vector(to_signed(-750,SDLEN)),
    to_std_logic_vector(to_signed(-772,SDLEN)),
    to_std_logic_vector(to_signed(-797,SDLEN)),
    to_std_logic_vector(to_signed(-827,SDLEN)),
    to_std_logic_vector(to_signed(-861,SDLEN)),
    to_std_logic_vector(to_signed(-901,SDLEN)),
    to_std_logic_vector(to_signed(-946,SDLEN)),
    to_std_logic_vector(to_signed(-998,SDLEN)),
    to_std_logic_vector(to_signed(-1059,SDLEN)),
    to_std_logic_vector(to_signed(-1132,SDLEN)),
    to_std_logic_vector(to_signed(-1219,SDLEN)),
    to_std_logic_vector(to_signed(-1322,SDLEN)),
    to_std_logic_vector(to_signed(-1450,SDLEN)),
    to_std_logic_vector(to_signed(-1608,SDLEN)),
    to_std_logic_vector(to_signed(-1811,SDLEN)),
    to_std_logic_vector(to_signed(-2081,SDLEN)),
    to_std_logic_vector(to_signed(-2444,SDLEN)),
    to_std_logic_vector(to_signed(-2979,SDLEN)),
    to_std_logic_vector(to_signed(-3813,SDLEN)),
    to_std_logic_vector(to_signed(-5323,SDLEN)),
    to_std_logic_vector(to_signed(-8812,SDLEN)),
    to_std_logic_vector(to_signed(-26887,SDLEN)),
    to_std_logic_vector(to_signed(32767,SDLEN)),
    to_std_logic_vector(to_signed(32729,SDLEN)),
    to_std_logic_vector(to_signed(32610,SDLEN)),
    to_std_logic_vector(to_signed(32413,SDLEN)),
    to_std_logic_vector(to_signed(32138,SDLEN)),
    to_std_logic_vector(to_signed(31786,SDLEN)),
    to_std_logic_vector(to_signed(31357,SDLEN)),
    to_std_logic_vector(to_signed(30853,SDLEN)),
    to_std_logic_vector(to_signed(30274,SDLEN)),
    to_std_logic_vector(to_signed(29622,SDLEN)),
    to_std_logic_vector(to_signed(28899,SDLEN)),
    to_std_logic_vector(to_signed(28106,SDLEN)),
    to_std_logic_vector(to_signed(27246,SDLEN)),
    to_std_logic_vector(to_signed(26320,SDLEN)),
    to_std_logic_vector(to_signed(25330,SDLEN)),
    to_std_logic_vector(to_signed(24279,SDLEN)),
    to_std_logic_vector(to_signed(23170,SDLEN)),
    to_std_logic_vector(to_signed(22006,SDLEN)),
    to_std_logic_vector(to_signed(20788,SDLEN)),
    to_std_logic_vector(to_signed(19520,SDLEN)),
    to_std_logic_vector(to_signed(18205,SDLEN)),
    to_std_logic_vector(to_signed(16846,SDLEN)),
    to_std_logic_vector(to_signed(15447,SDLEN)),
    to_std_logic_vector(to_signed(14010,SDLEN)),
    to_std_logic_vector(to_signed(12540,SDLEN)),
    to_std_logic_vector(to_signed(11039,SDLEN)),
    to_std_logic_vector(to_signed(9512,SDLEN)),
    to_std_logic_vector(to_signed(7962,SDLEN)),
    to_std_logic_vector(to_signed(6393,SDLEN)),
    to_std_logic_vector(to_signed(4808,SDLEN)),
    to_std_logic_vector(to_signed(3212,SDLEN)),
    to_std_logic_vector(to_signed(1608,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(-1608,SDLEN)),
    to_std_logic_vector(to_signed(-3212,SDLEN)),
    to_std_logic_vector(to_signed(-4808,SDLEN)),
    to_std_logic_vector(to_signed(-6393,SDLEN)),
    to_std_logic_vector(to_signed(-7962,SDLEN)),
    to_std_logic_vector(to_signed(-9512,SDLEN)),
    to_std_logic_vector(to_signed(-11039,SDLEN)),
    to_std_logic_vector(to_signed(-12540,SDLEN)),
    to_std_logic_vector(to_signed(-14010,SDLEN)),
    to_std_logic_vector(to_signed(-15447,SDLEN)),
    to_std_logic_vector(to_signed(-16846,SDLEN)),
    to_std_logic_vector(to_signed(-18205,SDLEN)),
    to_std_logic_vector(to_signed(-19520,SDLEN)),
    to_std_logic_vector(to_signed(-20788,SDLEN)),
    to_std_logic_vector(to_signed(-22006,SDLEN)),
    to_std_logic_vector(to_signed(-23170,SDLEN)),
    to_std_logic_vector(to_signed(-24279,SDLEN)),
    to_std_logic_vector(to_signed(-25330,SDLEN)),
    to_std_logic_vector(to_signed(-26320,SDLEN)),
    to_std_logic_vector(to_signed(-27246,SDLEN)),
    to_std_logic_vector(to_signed(-28106,SDLEN)),
    to_std_logic_vector(to_signed(-28899,SDLEN)),
    to_std_logic_vector(to_signed(-29622,SDLEN)),
    to_std_logic_vector(to_signed(-30274,SDLEN)),
    to_std_logic_vector(to_signed(-30853,SDLEN)),
    to_std_logic_vector(to_signed(-31357,SDLEN)),
    to_std_logic_vector(to_signed(-31786,SDLEN)),
    to_std_logic_vector(to_signed(-32138,SDLEN)),
    to_std_logic_vector(to_signed(-32413,SDLEN)),
    to_std_logic_vector(to_signed(-32610,SDLEN)),
    to_std_logic_vector(to_signed(-32729,SDLEN)),
    to_std_logic_vector(to_signed(-632,SDLEN)),
    to_std_logic_vector(to_signed(-1893,SDLEN)),
    to_std_logic_vector(to_signed(-3150,SDLEN)),
    to_std_logic_vector(to_signed(-4399,SDLEN)),
    to_std_logic_vector(to_signed(-5638,SDLEN)),
    to_std_logic_vector(to_signed(-6863,SDLEN)),
    to_std_logic_vector(to_signed(-8072,SDLEN)),
    to_std_logic_vector(to_signed(-9261,SDLEN)),
    to_std_logic_vector(to_signed(-10428,SDLEN)),
    to_std_logic_vector(to_signed(-11570,SDLEN)),
    to_std_logic_vector(to_signed(-12684,SDLEN)),
    to_std_logic_vector(to_signed(-13767,SDLEN)),
    to_std_logic_vector(to_signed(-14817,SDLEN)),
    to_std_logic_vector(to_signed(-15832,SDLEN)),
    to_std_logic_vector(to_signed(-16808,SDLEN)),
    to_std_logic_vector(to_signed(-17744,SDLEN)),
    to_std_logic_vector(to_signed(-18637,SDLEN)),
    to_std_logic_vector(to_signed(-19486,SDLEN)),
    to_std_logic_vector(to_signed(-20287,SDLEN)),
    to_std_logic_vector(to_signed(-21039,SDLEN)),
    to_std_logic_vector(to_signed(-21741,SDLEN)),
    to_std_logic_vector(to_signed(-22390,SDLEN)),
    to_std_logic_vector(to_signed(-22986,SDLEN)),
    to_std_logic_vector(to_signed(-23526,SDLEN)),
    to_std_logic_vector(to_signed(-24009,SDLEN)),
    to_std_logic_vector(to_signed(-24435,SDLEN)),
    to_std_logic_vector(to_signed(-24801,SDLEN)),
    to_std_logic_vector(to_signed(-25108,SDLEN)),
    to_std_logic_vector(to_signed(-25354,SDLEN)),
    to_std_logic_vector(to_signed(-25540,SDLEN)),
    to_std_logic_vector(to_signed(-25664,SDLEN)),
    to_std_logic_vector(to_signed(-25726,SDLEN)),
    to_std_logic_vector(to_signed(-25726,SDLEN)),
    to_std_logic_vector(to_signed(-25664,SDLEN)),
    to_std_logic_vector(to_signed(-25540,SDLEN)),
    to_std_logic_vector(to_signed(-25354,SDLEN)),
    to_std_logic_vector(to_signed(-25108,SDLEN)),
    to_std_logic_vector(to_signed(-24801,SDLEN)),
    to_std_logic_vector(to_signed(-24435,SDLEN)),
    to_std_logic_vector(to_signed(-24009,SDLEN)),
    to_std_logic_vector(to_signed(-23526,SDLEN)),
    to_std_logic_vector(to_signed(-22986,SDLEN)),
    to_std_logic_vector(to_signed(-22390,SDLEN)),
    to_std_logic_vector(to_signed(-21741,SDLEN)),
    to_std_logic_vector(to_signed(-21039,SDLEN)),
    to_std_logic_vector(to_signed(-20287,SDLEN)),
    to_std_logic_vector(to_signed(-19486,SDLEN)),
    to_std_logic_vector(to_signed(-18637,SDLEN)),
    to_std_logic_vector(to_signed(-17744,SDLEN)),
    to_std_logic_vector(to_signed(-16808,SDLEN)),
    to_std_logic_vector(to_signed(-15832,SDLEN)),
    to_std_logic_vector(to_signed(-14817,SDLEN)),
    to_std_logic_vector(to_signed(-13767,SDLEN)),
    to_std_logic_vector(to_signed(-12684,SDLEN)),
    to_std_logic_vector(to_signed(-11570,SDLEN)),
    to_std_logic_vector(to_signed(-10428,SDLEN)),
    to_std_logic_vector(to_signed(-9261,SDLEN)),
    to_std_logic_vector(to_signed(-8072,SDLEN)),
    to_std_logic_vector(to_signed(-6863,SDLEN)),
    to_std_logic_vector(to_signed(-5638,SDLEN)),
    to_std_logic_vector(to_signed(-4399,SDLEN)),
    to_std_logic_vector(to_signed(-3150,SDLEN)),
    to_std_logic_vector(to_signed(-1893,SDLEN)),
    to_std_logic_vector(to_signed(-632,SDLEN)),
    to_std_logic_vector(to_signed(-26887,SDLEN)),
    to_std_logic_vector(to_signed(-8812,SDLEN)),
    to_std_logic_vector(to_signed(-5323,SDLEN)),
    to_std_logic_vector(to_signed(-3813,SDLEN)),
    to_std_logic_vector(to_signed(-2979,SDLEN)),
    to_std_logic_vector(to_signed(-2444,SDLEN)),
    to_std_logic_vector(to_signed(-2081,SDLEN)),
    to_std_logic_vector(to_signed(-1811,SDLEN)),
    to_std_logic_vector(to_signed(-1608,SDLEN)),
    to_std_logic_vector(to_signed(-1450,SDLEN)),
    to_std_logic_vector(to_signed(-1322,SDLEN)),
    to_std_logic_vector(to_signed(-1219,SDLEN)),
    to_std_logic_vector(to_signed(-1132,SDLEN)),
    to_std_logic_vector(to_signed(-1059,SDLEN)),
    to_std_logic_vector(to_signed(-998,SDLEN)),
    to_std_logic_vector(to_signed(-946,SDLEN)),
    to_std_logic_vector(to_signed(-901,SDLEN)),
    to_std_logic_vector(to_signed(-861,SDLEN)),
    to_std_logic_vector(to_signed(-827,SDLEN)),
    to_std_logic_vector(to_signed(-797,SDLEN)),
    to_std_logic_vector(to_signed(-772,SDLEN)),
    to_std_logic_vector(to_signed(-750,SDLEN)),
    to_std_logic_vector(to_signed(-730,SDLEN)),
    to_std_logic_vector(to_signed(-713,SDLEN)),
    to_std_logic_vector(to_signed(-699,SDLEN)),
    to_std_logic_vector(to_signed(-687,SDLEN)),
    to_std_logic_vector(to_signed(-677,SDLEN)),
    to_std_logic_vector(to_signed(-668,SDLEN)),
    to_std_logic_vector(to_signed(-662,SDLEN)),
    to_std_logic_vector(to_signed(-657,SDLEN)),
    to_std_logic_vector(to_signed(-654,SDLEN)),
    to_std_logic_vector(to_signed(-652,SDLEN)),
    to_std_logic_vector(to_signed(-652,SDLEN)),
    to_std_logic_vector(to_signed(-654,SDLEN)),
    to_std_logic_vector(to_signed(-657,SDLEN)),
    to_std_logic_vector(to_signed(-662,SDLEN)),
    to_std_logic_vector(to_signed(-668,SDLEN)),
    to_std_logic_vector(to_signed(-677,SDLEN)),
    to_std_logic_vector(to_signed(-687,SDLEN)),
    to_std_logic_vector(to_signed(-699,SDLEN)),
    to_std_logic_vector(to_signed(-713,SDLEN)),
    to_std_logic_vector(to_signed(-730,SDLEN)),
    to_std_logic_vector(to_signed(-750,SDLEN)),
    to_std_logic_vector(to_signed(-772,SDLEN)),
    to_std_logic_vector(to_signed(-797,SDLEN)),
    to_std_logic_vector(to_signed(-827,SDLEN)),
    to_std_logic_vector(to_signed(-861,SDLEN)),
    to_std_logic_vector(to_signed(-901,SDLEN)),
    to_std_logic_vector(to_signed(-946,SDLEN)),
    to_std_logic_vector(to_signed(-998,SDLEN)),
    to_std_logic_vector(to_signed(-1059,SDLEN)),
    to_std_logic_vector(to_signed(-1132,SDLEN)),
    to_std_logic_vector(to_signed(-1219,SDLEN)),
    to_std_logic_vector(to_signed(-1322,SDLEN)),
    to_std_logic_vector(to_signed(-1450,SDLEN)),
    to_std_logic_vector(to_signed(-1608,SDLEN)),
    to_std_logic_vector(to_signed(-1811,SDLEN)),
    to_std_logic_vector(to_signed(-2081,SDLEN)),
    to_std_logic_vector(to_signed(-2444,SDLEN)),
    to_std_logic_vector(to_signed(-2979,SDLEN)),
    to_std_logic_vector(to_signed(-3813,SDLEN)),
    to_std_logic_vector(to_signed(-5323,SDLEN)),
    to_std_logic_vector(to_signed(-8812,SDLEN)),
    to_std_logic_vector(to_signed(-26887,SDLEN)),
    to_std_logic_vector(to_signed(1486,SDLEN)),
    to_std_logic_vector(to_signed(2168,SDLEN)),
    to_std_logic_vector(to_signed(3751,SDLEN)),
    to_std_logic_vector(to_signed(9074,SDLEN)),
    to_std_logic_vector(to_signed(12134,SDLEN)),
    to_std_logic_vector(to_signed(13944,SDLEN)),
    to_std_logic_vector(to_signed(17983,SDLEN)),
    to_std_logic_vector(to_signed(19173,SDLEN)),
    to_std_logic_vector(to_signed(21190,SDLEN)),
    to_std_logic_vector(to_signed(21820,SDLEN)),
    to_std_logic_vector(to_signed(1730,SDLEN)),
    to_std_logic_vector(to_signed(2640,SDLEN)),
    to_std_logic_vector(to_signed(3450,SDLEN)),
    to_std_logic_vector(to_signed(4870,SDLEN)),
    to_std_logic_vector(to_signed(6126,SDLEN)),
    to_std_logic_vector(to_signed(7876,SDLEN)),
    to_std_logic_vector(to_signed(15644,SDLEN)),
    to_std_logic_vector(to_signed(17817,SDLEN)),
    to_std_logic_vector(to_signed(20294,SDLEN)),
    to_std_logic_vector(to_signed(21902,SDLEN)),
    to_std_logic_vector(to_signed(1568,SDLEN)),
    to_std_logic_vector(to_signed(2256,SDLEN)),
    to_std_logic_vector(to_signed(3088,SDLEN)),
    to_std_logic_vector(to_signed(4874,SDLEN)),
    to_std_logic_vector(to_signed(11063,SDLEN)),
    to_std_logic_vector(to_signed(13393,SDLEN)),
    to_std_logic_vector(to_signed(18307,SDLEN)),
    to_std_logic_vector(to_signed(19293,SDLEN)),
    to_std_logic_vector(to_signed(21109,SDLEN)),
    to_std_logic_vector(to_signed(21741,SDLEN)),
    to_std_logic_vector(to_signed(1733,SDLEN)),
    to_std_logic_vector(to_signed(2512,SDLEN)),
    to_std_logic_vector(to_signed(3357,SDLEN)),
    to_std_logic_vector(to_signed(4708,SDLEN)),
    to_std_logic_vector(to_signed(6977,SDLEN)),
    to_std_logic_vector(to_signed(10296,SDLEN)),
    to_std_logic_vector(to_signed(17024,SDLEN)),
    to_std_logic_vector(to_signed(17956,SDLEN)),
    to_std_logic_vector(to_signed(19145,SDLEN)),
    to_std_logic_vector(to_signed(20350,SDLEN)),
    to_std_logic_vector(to_signed(1744,SDLEN)),
    to_std_logic_vector(to_signed(2436,SDLEN)),
    to_std_logic_vector(to_signed(3308,SDLEN)),
    to_std_logic_vector(to_signed(8731,SDLEN)),
    to_std_logic_vector(to_signed(10432,SDLEN)),
    to_std_logic_vector(to_signed(12007,SDLEN)),
    to_std_logic_vector(to_signed(15614,SDLEN)),
    to_std_logic_vector(to_signed(16639,SDLEN)),
    to_std_logic_vector(to_signed(21359,SDLEN)),
    to_std_logic_vector(to_signed(21913,SDLEN)),
    to_std_logic_vector(to_signed(1786,SDLEN)),
    to_std_logic_vector(to_signed(2369,SDLEN)),
    to_std_logic_vector(to_signed(3372,SDLEN)),
    to_std_logic_vector(to_signed(4521,SDLEN)),
    to_std_logic_vector(to_signed(6795,SDLEN)),
    to_std_logic_vector(to_signed(12963,SDLEN)),
    to_std_logic_vector(to_signed(17674,SDLEN)),
    to_std_logic_vector(to_signed(18988,SDLEN)),
    to_std_logic_vector(to_signed(20855,SDLEN)),
    to_std_logic_vector(to_signed(21640,SDLEN)),
    to_std_logic_vector(to_signed(1631,SDLEN)),
    to_std_logic_vector(to_signed(2433,SDLEN)),
    to_std_logic_vector(to_signed(3361,SDLEN)),
    to_std_logic_vector(to_signed(6328,SDLEN)),
    to_std_logic_vector(to_signed(10709,SDLEN)),
    to_std_logic_vector(to_signed(12013,SDLEN)),
    to_std_logic_vector(to_signed(13277,SDLEN)),
    to_std_logic_vector(to_signed(13904,SDLEN)),
    to_std_logic_vector(to_signed(19441,SDLEN)),
    to_std_logic_vector(to_signed(21088,SDLEN)),
    to_std_logic_vector(to_signed(1489,SDLEN)),
    to_std_logic_vector(to_signed(2364,SDLEN)),
    to_std_logic_vector(to_signed(3291,SDLEN)),
    to_std_logic_vector(to_signed(6250,SDLEN)),
    to_std_logic_vector(to_signed(9227,SDLEN)),
    to_std_logic_vector(to_signed(10403,SDLEN)),
    to_std_logic_vector(to_signed(13843,SDLEN)),
    to_std_logic_vector(to_signed(15278,SDLEN)),
    to_std_logic_vector(to_signed(17721,SDLEN)),
    to_std_logic_vector(to_signed(21451,SDLEN)),
    to_std_logic_vector(to_signed(1869,SDLEN)),
    to_std_logic_vector(to_signed(2533,SDLEN)),
    to_std_logic_vector(to_signed(3475,SDLEN)),
    to_std_logic_vector(to_signed(4365,SDLEN)),
    to_std_logic_vector(to_signed(9152,SDLEN)),
    to_std_logic_vector(to_signed(14513,SDLEN)),
    to_std_logic_vector(to_signed(15908,SDLEN)),
    to_std_logic_vector(to_signed(17022,SDLEN)),
    to_std_logic_vector(to_signed(20611,SDLEN)),
    to_std_logic_vector(to_signed(21411,SDLEN)),
    to_std_logic_vector(to_signed(2070,SDLEN)),
    to_std_logic_vector(to_signed(3025,SDLEN)),
    to_std_logic_vector(to_signed(4333,SDLEN)),
    to_std_logic_vector(to_signed(5854,SDLEN)),
    to_std_logic_vector(to_signed(7805,SDLEN)),
    to_std_logic_vector(to_signed(9231,SDLEN)),
    to_std_logic_vector(to_signed(10597,SDLEN)),
    to_std_logic_vector(to_signed(16047,SDLEN)),
    to_std_logic_vector(to_signed(20109,SDLEN)),
    to_std_logic_vector(to_signed(21834,SDLEN)),
    to_std_logic_vector(to_signed(1910,SDLEN)),
    to_std_logic_vector(to_signed(2673,SDLEN)),
    to_std_logic_vector(to_signed(3419,SDLEN)),
    to_std_logic_vector(to_signed(4261,SDLEN)),
    to_std_logic_vector(to_signed(11168,SDLEN)),
    to_std_logic_vector(to_signed(15111,SDLEN)),
    to_std_logic_vector(to_signed(16577,SDLEN)),
    to_std_logic_vector(to_signed(17591,SDLEN)),
    to_std_logic_vector(to_signed(19310,SDLEN)),
    to_std_logic_vector(to_signed(20265,SDLEN)),
    to_std_logic_vector(to_signed(1141,SDLEN)),
    to_std_logic_vector(to_signed(1815,SDLEN)),
    to_std_logic_vector(to_signed(2624,SDLEN)),
    to_std_logic_vector(to_signed(4623,SDLEN)),
    to_std_logic_vector(to_signed(6495,SDLEN)),
    to_std_logic_vector(to_signed(9588,SDLEN)),
    to_std_logic_vector(to_signed(13968,SDLEN)),
    to_std_logic_vector(to_signed(16428,SDLEN)),
    to_std_logic_vector(to_signed(19351,SDLEN)),
    to_std_logic_vector(to_signed(21286,SDLEN)),
    to_std_logic_vector(to_signed(2192,SDLEN)),
    to_std_logic_vector(to_signed(3171,SDLEN)),
    to_std_logic_vector(to_signed(4707,SDLEN)),
    to_std_logic_vector(to_signed(5808,SDLEN)),
    to_std_logic_vector(to_signed(10904,SDLEN)),
    to_std_logic_vector(to_signed(12500,SDLEN)),
    to_std_logic_vector(to_signed(14162,SDLEN)),
    to_std_logic_vector(to_signed(15664,SDLEN)),
    to_std_logic_vector(to_signed(21124,SDLEN)),
    to_std_logic_vector(to_signed(21789,SDLEN)),
    to_std_logic_vector(to_signed(1286,SDLEN)),
    to_std_logic_vector(to_signed(1907,SDLEN)),
    to_std_logic_vector(to_signed(2548,SDLEN)),
    to_std_logic_vector(to_signed(3453,SDLEN)),
    to_std_logic_vector(to_signed(9574,SDLEN)),
    to_std_logic_vector(to_signed(11964,SDLEN)),
    to_std_logic_vector(to_signed(15978,SDLEN)),
    to_std_logic_vector(to_signed(17344,SDLEN)),
    to_std_logic_vector(to_signed(19691,SDLEN)),
    to_std_logic_vector(to_signed(22495,SDLEN)),
    to_std_logic_vector(to_signed(1921,SDLEN)),
    to_std_logic_vector(to_signed(2720,SDLEN)),
    to_std_logic_vector(to_signed(4604,SDLEN)),
    to_std_logic_vector(to_signed(6684,SDLEN)),
    to_std_logic_vector(to_signed(11503,SDLEN)),
    to_std_logic_vector(to_signed(12992,SDLEN)),
    to_std_logic_vector(to_signed(14350,SDLEN)),
    to_std_logic_vector(to_signed(15262,SDLEN)),
    to_std_logic_vector(to_signed(16997,SDLEN)),
    to_std_logic_vector(to_signed(20791,SDLEN)),
    to_std_logic_vector(to_signed(2052,SDLEN)),
    to_std_logic_vector(to_signed(2759,SDLEN)),
    to_std_logic_vector(to_signed(3897,SDLEN)),
    to_std_logic_vector(to_signed(5246,SDLEN)),
    to_std_logic_vector(to_signed(6638,SDLEN)),
    to_std_logic_vector(to_signed(10267,SDLEN)),
    to_std_logic_vector(to_signed(15834,SDLEN)),
    to_std_logic_vector(to_signed(16814,SDLEN)),
    to_std_logic_vector(to_signed(18149,SDLEN)),
    to_std_logic_vector(to_signed(21675,SDLEN)),
    to_std_logic_vector(to_signed(1798,SDLEN)),
    to_std_logic_vector(to_signed(2497,SDLEN)),
    to_std_logic_vector(to_signed(5617,SDLEN)),
    to_std_logic_vector(to_signed(11449,SDLEN)),
    to_std_logic_vector(to_signed(13189,SDLEN)),
    to_std_logic_vector(to_signed(14711,SDLEN)),
    to_std_logic_vector(to_signed(17050,SDLEN)),
    to_std_logic_vector(to_signed(18195,SDLEN)),
    to_std_logic_vector(to_signed(20307,SDLEN)),
    to_std_logic_vector(to_signed(21182,SDLEN)),
    to_std_logic_vector(to_signed(1009,SDLEN)),
    to_std_logic_vector(to_signed(1647,SDLEN)),
    to_std_logic_vector(to_signed(2889,SDLEN)),
    to_std_logic_vector(to_signed(5709,SDLEN)),
    to_std_logic_vector(to_signed(9541,SDLEN)),
    to_std_logic_vector(to_signed(12354,SDLEN)),
    to_std_logic_vector(to_signed(15231,SDLEN)),
    to_std_logic_vector(to_signed(18494,SDLEN)),
    to_std_logic_vector(to_signed(20966,SDLEN)),
    to_std_logic_vector(to_signed(22033,SDLEN)),
    to_std_logic_vector(to_signed(3016,SDLEN)),
    to_std_logic_vector(to_signed(3794,SDLEN)),
    to_std_logic_vector(to_signed(5406,SDLEN)),
    to_std_logic_vector(to_signed(7469,SDLEN)),
    to_std_logic_vector(to_signed(12488,SDLEN)),
    to_std_logic_vector(to_signed(13984,SDLEN)),
    to_std_logic_vector(to_signed(15328,SDLEN)),
    to_std_logic_vector(to_signed(16334,SDLEN)),
    to_std_logic_vector(to_signed(19952,SDLEN)),
    to_std_logic_vector(to_signed(20791,SDLEN)),
    to_std_logic_vector(to_signed(2203,SDLEN)),
    to_std_logic_vector(to_signed(3040,SDLEN)),
    to_std_logic_vector(to_signed(3796,SDLEN)),
    to_std_logic_vector(to_signed(5442,SDLEN)),
    to_std_logic_vector(to_signed(11987,SDLEN)),
    to_std_logic_vector(to_signed(13512,SDLEN)),
    to_std_logic_vector(to_signed(14931,SDLEN)),
    to_std_logic_vector(to_signed(16370,SDLEN)),
    to_std_logic_vector(to_signed(17856,SDLEN)),
    to_std_logic_vector(to_signed(18803,SDLEN)),
    to_std_logic_vector(to_signed(2912,SDLEN)),
    to_std_logic_vector(to_signed(4292,SDLEN)),
    to_std_logic_vector(to_signed(7988,SDLEN)),
    to_std_logic_vector(to_signed(9572,SDLEN)),
    to_std_logic_vector(to_signed(11562,SDLEN)),
    to_std_logic_vector(to_signed(13244,SDLEN)),
    to_std_logic_vector(to_signed(14556,SDLEN)),
    to_std_logic_vector(to_signed(16529,SDLEN)),
    to_std_logic_vector(to_signed(20004,SDLEN)),
    to_std_logic_vector(to_signed(21073,SDLEN)),
    to_std_logic_vector(to_signed(2861,SDLEN)),
    to_std_logic_vector(to_signed(3607,SDLEN)),
    to_std_logic_vector(to_signed(5923,SDLEN)),
    to_std_logic_vector(to_signed(7034,SDLEN)),
    to_std_logic_vector(to_signed(9234,SDLEN)),
    to_std_logic_vector(to_signed(12054,SDLEN)),
    to_std_logic_vector(to_signed(13729,SDLEN)),
    to_std_logic_vector(to_signed(18056,SDLEN)),
    to_std_logic_vector(to_signed(20262,SDLEN)),
    to_std_logic_vector(to_signed(20974,SDLEN)),
    to_std_logic_vector(to_signed(3069,SDLEN)),
    to_std_logic_vector(to_signed(4311,SDLEN)),
    to_std_logic_vector(to_signed(5967,SDLEN)),
    to_std_logic_vector(to_signed(7367,SDLEN)),
    to_std_logic_vector(to_signed(11482,SDLEN)),
    to_std_logic_vector(to_signed(12699,SDLEN)),
    to_std_logic_vector(to_signed(14309,SDLEN)),
    to_std_logic_vector(to_signed(16233,SDLEN)),
    to_std_logic_vector(to_signed(18333,SDLEN)),
    to_std_logic_vector(to_signed(19172,SDLEN)),
    to_std_logic_vector(to_signed(2434,SDLEN)),
    to_std_logic_vector(to_signed(3661,SDLEN)),
    to_std_logic_vector(to_signed(4866,SDLEN)),
    to_std_logic_vector(to_signed(5798,SDLEN)),
    to_std_logic_vector(to_signed(10383,SDLEN)),
    to_std_logic_vector(to_signed(11722,SDLEN)),
    to_std_logic_vector(to_signed(13049,SDLEN)),
    to_std_logic_vector(to_signed(15668,SDLEN)),
    to_std_logic_vector(to_signed(18862,SDLEN)),
    to_std_logic_vector(to_signed(19831,SDLEN)),
    to_std_logic_vector(to_signed(2020,SDLEN)),
    to_std_logic_vector(to_signed(2605,SDLEN)),
    to_std_logic_vector(to_signed(3860,SDLEN)),
    to_std_logic_vector(to_signed(9241,SDLEN)),
    to_std_logic_vector(to_signed(13275,SDLEN)),
    to_std_logic_vector(to_signed(14644,SDLEN)),
    to_std_logic_vector(to_signed(16010,SDLEN)),
    to_std_logic_vector(to_signed(17099,SDLEN)),
    to_std_logic_vector(to_signed(19268,SDLEN)),
    to_std_logic_vector(to_signed(20251,SDLEN)),
    to_std_logic_vector(to_signed(1877,SDLEN)),
    to_std_logic_vector(to_signed(2809,SDLEN)),
    to_std_logic_vector(to_signed(3590,SDLEN)),
    to_std_logic_vector(to_signed(4707,SDLEN)),
    to_std_logic_vector(to_signed(11056,SDLEN)),
    to_std_logic_vector(to_signed(12441,SDLEN)),
    to_std_logic_vector(to_signed(15622,SDLEN)),
    to_std_logic_vector(to_signed(17168,SDLEN)),
    to_std_logic_vector(to_signed(18761,SDLEN)),
    to_std_logic_vector(to_signed(19907,SDLEN)),
    to_std_logic_vector(to_signed(2107,SDLEN)),
    to_std_logic_vector(to_signed(2873,SDLEN)),
    to_std_logic_vector(to_signed(3673,SDLEN)),
    to_std_logic_vector(to_signed(5799,SDLEN)),
    to_std_logic_vector(to_signed(13579,SDLEN)),
    to_std_logic_vector(to_signed(14687,SDLEN)),
    to_std_logic_vector(to_signed(15938,SDLEN)),
    to_std_logic_vector(to_signed(17077,SDLEN)),
    to_std_logic_vector(to_signed(18890,SDLEN)),
    to_std_logic_vector(to_signed(19831,SDLEN)),
    to_std_logic_vector(to_signed(1612,SDLEN)),
    to_std_logic_vector(to_signed(2284,SDLEN)),
    to_std_logic_vector(to_signed(2944,SDLEN)),
    to_std_logic_vector(to_signed(3572,SDLEN)),
    to_std_logic_vector(to_signed(8219,SDLEN)),
    to_std_logic_vector(to_signed(13959,SDLEN)),
    to_std_logic_vector(to_signed(15924,SDLEN)),
    to_std_logic_vector(to_signed(17239,SDLEN)),
    to_std_logic_vector(to_signed(18592,SDLEN)),
    to_std_logic_vector(to_signed(20117,SDLEN)),
    to_std_logic_vector(to_signed(2420,SDLEN)),
    to_std_logic_vector(to_signed(3156,SDLEN)),
    to_std_logic_vector(to_signed(6542,SDLEN)),
    to_std_logic_vector(to_signed(10215,SDLEN)),
    to_std_logic_vector(to_signed(12061,SDLEN)),
    to_std_logic_vector(to_signed(13534,SDLEN)),
    to_std_logic_vector(to_signed(15305,SDLEN)),
    to_std_logic_vector(to_signed(16452,SDLEN)),
    to_std_logic_vector(to_signed(18717,SDLEN)),
    to_std_logic_vector(to_signed(19880,SDLEN)),
    to_std_logic_vector(to_signed(1667,SDLEN)),
    to_std_logic_vector(to_signed(2612,SDLEN)),
    to_std_logic_vector(to_signed(3534,SDLEN)),
    to_std_logic_vector(to_signed(5237,SDLEN)),
    to_std_logic_vector(to_signed(10513,SDLEN)),
    to_std_logic_vector(to_signed(11696,SDLEN)),
    to_std_logic_vector(to_signed(12940,SDLEN)),
    to_std_logic_vector(to_signed(16798,SDLEN)),
    to_std_logic_vector(to_signed(18058,SDLEN)),
    to_std_logic_vector(to_signed(19378,SDLEN)),
    to_std_logic_vector(to_signed(2388,SDLEN)),
    to_std_logic_vector(to_signed(3017,SDLEN)),
    to_std_logic_vector(to_signed(4839,SDLEN)),
    to_std_logic_vector(to_signed(9333,SDLEN)),
    to_std_logic_vector(to_signed(11413,SDLEN)),
    to_std_logic_vector(to_signed(12730,SDLEN)),
    to_std_logic_vector(to_signed(15024,SDLEN)),
    to_std_logic_vector(to_signed(16248,SDLEN)),
    to_std_logic_vector(to_signed(17449,SDLEN)),
    to_std_logic_vector(to_signed(18677,SDLEN)),
    to_std_logic_vector(to_signed(1875,SDLEN)),
    to_std_logic_vector(to_signed(2786,SDLEN)),
    to_std_logic_vector(to_signed(4231,SDLEN)),
    to_std_logic_vector(to_signed(6320,SDLEN)),
    to_std_logic_vector(to_signed(8694,SDLEN)),
    to_std_logic_vector(to_signed(10149,SDLEN)),
    to_std_logic_vector(to_signed(11785,SDLEN)),
    to_std_logic_vector(to_signed(17013,SDLEN)),
    to_std_logic_vector(to_signed(18608,SDLEN)),
    to_std_logic_vector(to_signed(19960,SDLEN)),
    to_std_logic_vector(to_signed(679,SDLEN)),
    to_std_logic_vector(to_signed(1411,SDLEN)),
    to_std_logic_vector(to_signed(4654,SDLEN)),
    to_std_logic_vector(to_signed(8006,SDLEN)),
    to_std_logic_vector(to_signed(11446,SDLEN)),
    to_std_logic_vector(to_signed(13249,SDLEN)),
    to_std_logic_vector(to_signed(15763,SDLEN)),
    to_std_logic_vector(to_signed(18127,SDLEN)),
    to_std_logic_vector(to_signed(20361,SDLEN)),
    to_std_logic_vector(to_signed(21567,SDLEN)),
    to_std_logic_vector(to_signed(1838,SDLEN)),
    to_std_logic_vector(to_signed(2596,SDLEN)),
    to_std_logic_vector(to_signed(3578,SDLEN)),
    to_std_logic_vector(to_signed(4608,SDLEN)),
    to_std_logic_vector(to_signed(5650,SDLEN)),
    to_std_logic_vector(to_signed(11274,SDLEN)),
    to_std_logic_vector(to_signed(14355,SDLEN)),
    to_std_logic_vector(to_signed(15886,SDLEN)),
    to_std_logic_vector(to_signed(20579,SDLEN)),
    to_std_logic_vector(to_signed(21754,SDLEN)),
    to_std_logic_vector(to_signed(1303,SDLEN)),
    to_std_logic_vector(to_signed(1955,SDLEN)),
    to_std_logic_vector(to_signed(2395,SDLEN)),
    to_std_logic_vector(to_signed(3322,SDLEN)),
    to_std_logic_vector(to_signed(12023,SDLEN)),
    to_std_logic_vector(to_signed(13764,SDLEN)),
    to_std_logic_vector(to_signed(15883,SDLEN)),
    to_std_logic_vector(to_signed(18077,SDLEN)),
    to_std_logic_vector(to_signed(20180,SDLEN)),
    to_std_logic_vector(to_signed(21232,SDLEN)),
    to_std_logic_vector(to_signed(1438,SDLEN)),
    to_std_logic_vector(to_signed(2102,SDLEN)),
    to_std_logic_vector(to_signed(2663,SDLEN)),
    to_std_logic_vector(to_signed(3462,SDLEN)),
    to_std_logic_vector(to_signed(8328,SDLEN)),
    to_std_logic_vector(to_signed(10362,SDLEN)),
    to_std_logic_vector(to_signed(13763,SDLEN)),
    to_std_logic_vector(to_signed(17248,SDLEN)),
    to_std_logic_vector(to_signed(19732,SDLEN)),
    to_std_logic_vector(to_signed(22344,SDLEN)),
    to_std_logic_vector(to_signed(860,SDLEN)),
    to_std_logic_vector(to_signed(1904,SDLEN)),
    to_std_logic_vector(to_signed(6098,SDLEN)),
    to_std_logic_vector(to_signed(7775,SDLEN)),
    to_std_logic_vector(to_signed(9815,SDLEN)),
    to_std_logic_vector(to_signed(12007,SDLEN)),
    to_std_logic_vector(to_signed(14821,SDLEN)),
    to_std_logic_vector(to_signed(16709,SDLEN)),
    to_std_logic_vector(to_signed(19787,SDLEN)),
    to_std_logic_vector(to_signed(21132,SDLEN)),
    to_std_logic_vector(to_signed(1673,SDLEN)),
    to_std_logic_vector(to_signed(2723,SDLEN)),
    to_std_logic_vector(to_signed(3704,SDLEN)),
    to_std_logic_vector(to_signed(6125,SDLEN)),
    to_std_logic_vector(to_signed(7668,SDLEN)),
    to_std_logic_vector(to_signed(9447,SDLEN)),
    to_std_logic_vector(to_signed(13683,SDLEN)),
    to_std_logic_vector(to_signed(14443,SDLEN)),
    to_std_logic_vector(to_signed(20538,SDLEN)),
    to_std_logic_vector(to_signed(21731,SDLEN)),
    to_std_logic_vector(to_signed(1246,SDLEN)),
    to_std_logic_vector(to_signed(1849,SDLEN)),
    to_std_logic_vector(to_signed(2902,SDLEN)),
    to_std_logic_vector(to_signed(4508,SDLEN)),
    to_std_logic_vector(to_signed(7221,SDLEN)),
    to_std_logic_vector(to_signed(12710,SDLEN)),
    to_std_logic_vector(to_signed(14835,SDLEN)),
    to_std_logic_vector(to_signed(16314,SDLEN)),
    to_std_logic_vector(to_signed(19335,SDLEN)),
    to_std_logic_vector(to_signed(22720,SDLEN)),
    to_std_logic_vector(to_signed(1525,SDLEN)),
    to_std_logic_vector(to_signed(2260,SDLEN)),
    to_std_logic_vector(to_signed(3862,SDLEN)),
    to_std_logic_vector(to_signed(5659,SDLEN)),
    to_std_logic_vector(to_signed(7342,SDLEN)),
    to_std_logic_vector(to_signed(11748,SDLEN)),
    to_std_logic_vector(to_signed(13370,SDLEN)),
    to_std_logic_vector(to_signed(14442,SDLEN)),
    to_std_logic_vector(to_signed(18044,SDLEN)),
    to_std_logic_vector(to_signed(21334,SDLEN)),
    to_std_logic_vector(to_signed(1196,SDLEN)),
    to_std_logic_vector(to_signed(1846,SDLEN)),
    to_std_logic_vector(to_signed(3104,SDLEN)),
    to_std_logic_vector(to_signed(7063,SDLEN)),
    to_std_logic_vector(to_signed(10972,SDLEN)),
    to_std_logic_vector(to_signed(12905,SDLEN)),
    to_std_logic_vector(to_signed(14814,SDLEN)),
    to_std_logic_vector(to_signed(17037,SDLEN)),
    to_std_logic_vector(to_signed(19922,SDLEN)),
    to_std_logic_vector(to_signed(22636,SDLEN)),
    to_std_logic_vector(to_signed(2147,SDLEN)),
    to_std_logic_vector(to_signed(3106,SDLEN)),
    to_std_logic_vector(to_signed(4475,SDLEN)),
    to_std_logic_vector(to_signed(6511,SDLEN)),
    to_std_logic_vector(to_signed(8227,SDLEN)),
    to_std_logic_vector(to_signed(9765,SDLEN)),
    to_std_logic_vector(to_signed(10984,SDLEN)),
    to_std_logic_vector(to_signed(12161,SDLEN)),
    to_std_logic_vector(to_signed(18971,SDLEN)),
    to_std_logic_vector(to_signed(21300,SDLEN)),
    to_std_logic_vector(to_signed(1585,SDLEN)),
    to_std_logic_vector(to_signed(2405,SDLEN)),
    to_std_logic_vector(to_signed(2994,SDLEN)),
    to_std_logic_vector(to_signed(4036,SDLEN)),
    to_std_logic_vector(to_signed(11481,SDLEN)),
    to_std_logic_vector(to_signed(13177,SDLEN)),
    to_std_logic_vector(to_signed(14519,SDLEN)),
    to_std_logic_vector(to_signed(15431,SDLEN)),
    to_std_logic_vector(to_signed(19967,SDLEN)),
    to_std_logic_vector(to_signed(21275,SDLEN)),
    to_std_logic_vector(to_signed(1778,SDLEN)),
    to_std_logic_vector(to_signed(2688,SDLEN)),
    to_std_logic_vector(to_signed(3614,SDLEN)),
    to_std_logic_vector(to_signed(4680,SDLEN)),
    to_std_logic_vector(to_signed(9465,SDLEN)),
    to_std_logic_vector(to_signed(11064,SDLEN)),
    to_std_logic_vector(to_signed(12473,SDLEN)),
    to_std_logic_vector(to_signed(16320,SDLEN)),
    to_std_logic_vector(to_signed(19742,SDLEN)),
    to_std_logic_vector(to_signed(20800,SDLEN)),
    to_std_logic_vector(to_signed(1862,SDLEN)),
    to_std_logic_vector(to_signed(2586,SDLEN)),
    to_std_logic_vector(to_signed(3492,SDLEN)),
    to_std_logic_vector(to_signed(6719,SDLEN)),
    to_std_logic_vector(to_signed(11708,SDLEN)),
    to_std_logic_vector(to_signed(13012,SDLEN)),
    to_std_logic_vector(to_signed(14364,SDLEN)),
    to_std_logic_vector(to_signed(16128,SDLEN)),
    to_std_logic_vector(to_signed(19610,SDLEN)),
    to_std_logic_vector(to_signed(20425,SDLEN)),
    to_std_logic_vector(to_signed(1395,SDLEN)),
    to_std_logic_vector(to_signed(2156,SDLEN)),
    to_std_logic_vector(to_signed(2669,SDLEN)),
    to_std_logic_vector(to_signed(3386,SDLEN)),
    to_std_logic_vector(to_signed(10607,SDLEN)),
    to_std_logic_vector(to_signed(12125,SDLEN)),
    to_std_logic_vector(to_signed(13614,SDLEN)),
    to_std_logic_vector(to_signed(16705,SDLEN)),
    to_std_logic_vector(to_signed(18976,SDLEN)),
    to_std_logic_vector(to_signed(21367,SDLEN)),
    to_std_logic_vector(to_signed(1444,SDLEN)),
    to_std_logic_vector(to_signed(2117,SDLEN)),
    to_std_logic_vector(to_signed(3286,SDLEN)),
    to_std_logic_vector(to_signed(6233,SDLEN)),
    to_std_logic_vector(to_signed(9423,SDLEN)),
    to_std_logic_vector(to_signed(12981,SDLEN)),
    to_std_logic_vector(to_signed(14998,SDLEN)),
    to_std_logic_vector(to_signed(15853,SDLEN)),
    to_std_logic_vector(to_signed(17188,SDLEN)),
    to_std_logic_vector(to_signed(21857,SDLEN)),
    to_std_logic_vector(to_signed(2004,SDLEN)),
    to_std_logic_vector(to_signed(2895,SDLEN)),
    to_std_logic_vector(to_signed(3783,SDLEN)),
    to_std_logic_vector(to_signed(4897,SDLEN)),
    to_std_logic_vector(to_signed(6168,SDLEN)),
    to_std_logic_vector(to_signed(7297,SDLEN)),
    to_std_logic_vector(to_signed(12609,SDLEN)),
    to_std_logic_vector(to_signed(16445,SDLEN)),
    to_std_logic_vector(to_signed(19297,SDLEN)),
    to_std_logic_vector(to_signed(21465,SDLEN)),
    to_std_logic_vector(to_signed(1495,SDLEN)),
    to_std_logic_vector(to_signed(2863,SDLEN)),
    to_std_logic_vector(to_signed(6360,SDLEN)),
    to_std_logic_vector(to_signed(8100,SDLEN)),
    to_std_logic_vector(to_signed(11399,SDLEN)),
    to_std_logic_vector(to_signed(14271,SDLEN)),
    to_std_logic_vector(to_signed(15902,SDLEN)),
    to_std_logic_vector(to_signed(17711,SDLEN)),
    to_std_logic_vector(to_signed(20479,SDLEN)),
    to_std_logic_vector(to_signed(22061,SDLEN)),
    to_std_logic_vector(to_signed(2484,SDLEN)),
    to_std_logic_vector(to_signed(3114,SDLEN)),
    to_std_logic_vector(to_signed(5718,SDLEN)),
    to_std_logic_vector(to_signed(7097,SDLEN)),
    to_std_logic_vector(to_signed(8400,SDLEN)),
    to_std_logic_vector(to_signed(12616,SDLEN)),
    to_std_logic_vector(to_signed(14073,SDLEN)),
    to_std_logic_vector(to_signed(14847,SDLEN)),
    to_std_logic_vector(to_signed(20535,SDLEN)),
    to_std_logic_vector(to_signed(21396,SDLEN)),
    to_std_logic_vector(to_signed(2424,SDLEN)),
    to_std_logic_vector(to_signed(3277,SDLEN)),
    to_std_logic_vector(to_signed(5296,SDLEN)),
    to_std_logic_vector(to_signed(6284,SDLEN)),
    to_std_logic_vector(to_signed(11290,SDLEN)),
    to_std_logic_vector(to_signed(12903,SDLEN)),
    to_std_logic_vector(to_signed(16022,SDLEN)),
    to_std_logic_vector(to_signed(17508,SDLEN)),
    to_std_logic_vector(to_signed(19333,SDLEN)),
    to_std_logic_vector(to_signed(20283,SDLEN)),
    to_std_logic_vector(to_signed(2565,SDLEN)),
    to_std_logic_vector(to_signed(3778,SDLEN)),
    to_std_logic_vector(to_signed(5360,SDLEN)),
    to_std_logic_vector(to_signed(6989,SDLEN)),
    to_std_logic_vector(to_signed(8782,SDLEN)),
    to_std_logic_vector(to_signed(10428,SDLEN)),
    to_std_logic_vector(to_signed(14390,SDLEN)),
    to_std_logic_vector(to_signed(15742,SDLEN)),
    to_std_logic_vector(to_signed(17770,SDLEN)),
    to_std_logic_vector(to_signed(21734,SDLEN)),
    to_std_logic_vector(to_signed(2727,SDLEN)),
    to_std_logic_vector(to_signed(3384,SDLEN)),
    to_std_logic_vector(to_signed(6613,SDLEN)),
    to_std_logic_vector(to_signed(9254,SDLEN)),
    to_std_logic_vector(to_signed(10542,SDLEN)),
    to_std_logic_vector(to_signed(12236,SDLEN)),
    to_std_logic_vector(to_signed(14651,SDLEN)),
    to_std_logic_vector(to_signed(15687,SDLEN)),
    to_std_logic_vector(to_signed(20074,SDLEN)),
    to_std_logic_vector(to_signed(21102,SDLEN)),
    to_std_logic_vector(to_signed(1916,SDLEN)),
    to_std_logic_vector(to_signed(2953,SDLEN)),
    to_std_logic_vector(to_signed(6274,SDLEN)),
    to_std_logic_vector(to_signed(8088,SDLEN)),
    to_std_logic_vector(to_signed(9710,SDLEN)),
    to_std_logic_vector(to_signed(10925,SDLEN)),
    to_std_logic_vector(to_signed(12392,SDLEN)),
    to_std_logic_vector(to_signed(16434,SDLEN)),
    to_std_logic_vector(to_signed(20010,SDLEN)),
    to_std_logic_vector(to_signed(21183,SDLEN)),
    to_std_logic_vector(to_signed(3384,SDLEN)),
    to_std_logic_vector(to_signed(4366,SDLEN)),
    to_std_logic_vector(to_signed(5349,SDLEN)),
    to_std_logic_vector(to_signed(7667,SDLEN)),
    to_std_logic_vector(to_signed(11180,SDLEN)),
    to_std_logic_vector(to_signed(12605,SDLEN)),
    to_std_logic_vector(to_signed(13921,SDLEN)),
    to_std_logic_vector(to_signed(15324,SDLEN)),
    to_std_logic_vector(to_signed(19901,SDLEN)),
    to_std_logic_vector(to_signed(20754,SDLEN)),
    to_std_logic_vector(to_signed(3075,SDLEN)),
    to_std_logic_vector(to_signed(4283,SDLEN)),
    to_std_logic_vector(to_signed(5951,SDLEN)),
    to_std_logic_vector(to_signed(7619,SDLEN)),
    to_std_logic_vector(to_signed(9604,SDLEN)),
    to_std_logic_vector(to_signed(11010,SDLEN)),
    to_std_logic_vector(to_signed(12384,SDLEN)),
    to_std_logic_vector(to_signed(14006,SDLEN)),
    to_std_logic_vector(to_signed(20658,SDLEN)),
    to_std_logic_vector(to_signed(21497,SDLEN)),
    to_std_logic_vector(to_signed(1751,SDLEN)),
    to_std_logic_vector(to_signed(2455,SDLEN)),
    to_std_logic_vector(to_signed(5147,SDLEN)),
    to_std_logic_vector(to_signed(9966,SDLEN)),
    to_std_logic_vector(to_signed(11621,SDLEN)),
    to_std_logic_vector(to_signed(13176,SDLEN)),
    to_std_logic_vector(to_signed(14739,SDLEN)),
    to_std_logic_vector(to_signed(16470,SDLEN)),
    to_std_logic_vector(to_signed(20788,SDLEN)),
    to_std_logic_vector(to_signed(21756,SDLEN)),
    to_std_logic_vector(to_signed(1442,SDLEN)),
    to_std_logic_vector(to_signed(2188,SDLEN)),
    to_std_logic_vector(to_signed(3330,SDLEN)),
    to_std_logic_vector(to_signed(6813,SDLEN)),
    to_std_logic_vector(to_signed(8929,SDLEN)),
    to_std_logic_vector(to_signed(12135,SDLEN)),
    to_std_logic_vector(to_signed(14476,SDLEN)),
    to_std_logic_vector(to_signed(15306,SDLEN)),
    to_std_logic_vector(to_signed(19635,SDLEN)),
    to_std_logic_vector(to_signed(20544,SDLEN)),
    to_std_logic_vector(to_signed(2294,SDLEN)),
    to_std_logic_vector(to_signed(2895,SDLEN)),
    to_std_logic_vector(to_signed(4070,SDLEN)),
    to_std_logic_vector(to_signed(8035,SDLEN)),
    to_std_logic_vector(to_signed(12233,SDLEN)),
    to_std_logic_vector(to_signed(13416,SDLEN)),
    to_std_logic_vector(to_signed(14762,SDLEN)),
    to_std_logic_vector(to_signed(17367,SDLEN)),
    to_std_logic_vector(to_signed(18952,SDLEN)),
    to_std_logic_vector(to_signed(19688,SDLEN)),
    to_std_logic_vector(to_signed(1937,SDLEN)),
    to_std_logic_vector(to_signed(2659,SDLEN)),
    to_std_logic_vector(to_signed(4602,SDLEN)),
    to_std_logic_vector(to_signed(6697,SDLEN)),
    to_std_logic_vector(to_signed(9071,SDLEN)),
    to_std_logic_vector(to_signed(12863,SDLEN)),
    to_std_logic_vector(to_signed(14197,SDLEN)),
    to_std_logic_vector(to_signed(15230,SDLEN)),
    to_std_logic_vector(to_signed(16047,SDLEN)),
    to_std_logic_vector(to_signed(18877,SDLEN)),
    to_std_logic_vector(to_signed(2071,SDLEN)),
    to_std_logic_vector(to_signed(2663,SDLEN)),
    to_std_logic_vector(to_signed(4216,SDLEN)),
    to_std_logic_vector(to_signed(9445,SDLEN)),
    to_std_logic_vector(to_signed(10887,SDLEN)),
    to_std_logic_vector(to_signed(12292,SDLEN)),
    to_std_logic_vector(to_signed(13949,SDLEN)),
    to_std_logic_vector(to_signed(14909,SDLEN)),
    to_std_logic_vector(to_signed(19236,SDLEN)),
    to_std_logic_vector(to_signed(20341,SDLEN)),
    to_std_logic_vector(to_signed(1740,SDLEN)),
    to_std_logic_vector(to_signed(2491,SDLEN)),
    to_std_logic_vector(to_signed(3488,SDLEN)),
    to_std_logic_vector(to_signed(8138,SDLEN)),
    to_std_logic_vector(to_signed(9656,SDLEN)),
    to_std_logic_vector(to_signed(11153,SDLEN)),
    to_std_logic_vector(to_signed(13206,SDLEN)),
    to_std_logic_vector(to_signed(14688,SDLEN)),
    to_std_logic_vector(to_signed(20896,SDLEN)),
    to_std_logic_vector(to_signed(21907,SDLEN)),
    to_std_logic_vector(to_signed(2199,SDLEN)),
    to_std_logic_vector(to_signed(2881,SDLEN)),
    to_std_logic_vector(to_signed(4675,SDLEN)),
    to_std_logic_vector(to_signed(8527,SDLEN)),
    to_std_logic_vector(to_signed(10051,SDLEN)),
    to_std_logic_vector(to_signed(11408,SDLEN)),
    to_std_logic_vector(to_signed(14435,SDLEN)),
    to_std_logic_vector(to_signed(15463,SDLEN)),
    to_std_logic_vector(to_signed(17190,SDLEN)),
    to_std_logic_vector(to_signed(20597,SDLEN)),
    to_std_logic_vector(to_signed(1943,SDLEN)),
    to_std_logic_vector(to_signed(2988,SDLEN)),
    to_std_logic_vector(to_signed(4177,SDLEN)),
    to_std_logic_vector(to_signed(6039,SDLEN)),
    to_std_logic_vector(to_signed(7478,SDLEN)),
    to_std_logic_vector(to_signed(8536,SDLEN)),
    to_std_logic_vector(to_signed(14181,SDLEN)),
    to_std_logic_vector(to_signed(15551,SDLEN)),
    to_std_logic_vector(to_signed(17622,SDLEN)),
    to_std_logic_vector(to_signed(21579,SDLEN)),
    to_std_logic_vector(to_signed(1825,SDLEN)),
    to_std_logic_vector(to_signed(3175,SDLEN)),
    to_std_logic_vector(to_signed(7062,SDLEN)),
    to_std_logic_vector(to_signed(9818,SDLEN)),
    to_std_logic_vector(to_signed(12824,SDLEN)),
    to_std_logic_vector(to_signed(15450,SDLEN)),
    to_std_logic_vector(to_signed(18330,SDLEN)),
    to_std_logic_vector(to_signed(19856,SDLEN)),
    to_std_logic_vector(to_signed(21830,SDLEN)),
    to_std_logic_vector(to_signed(22412,SDLEN)),
    to_std_logic_vector(to_signed(2464,SDLEN)),
    to_std_logic_vector(to_signed(3046,SDLEN)),
    to_std_logic_vector(to_signed(4822,SDLEN)),
    to_std_logic_vector(to_signed(5977,SDLEN)),
    to_std_logic_vector(to_signed(7696,SDLEN)),
    to_std_logic_vector(to_signed(15398,SDLEN)),
    to_std_logic_vector(to_signed(16730,SDLEN)),
    to_std_logic_vector(to_signed(17646,SDLEN)),
    to_std_logic_vector(to_signed(20588,SDLEN)),
    to_std_logic_vector(to_signed(21320,SDLEN)),
    to_std_logic_vector(to_signed(2550,SDLEN)),
    to_std_logic_vector(to_signed(3393,SDLEN)),
    to_std_logic_vector(to_signed(5305,SDLEN)),
    to_std_logic_vector(to_signed(6920,SDLEN)),
    to_std_logic_vector(to_signed(10235,SDLEN)),
    to_std_logic_vector(to_signed(14083,SDLEN)),
    to_std_logic_vector(to_signed(18143,SDLEN)),
    to_std_logic_vector(to_signed(19195,SDLEN)),
    to_std_logic_vector(to_signed(20681,SDLEN)),
    to_std_logic_vector(to_signed(21336,SDLEN)),
    to_std_logic_vector(to_signed(3003,SDLEN)),
    to_std_logic_vector(to_signed(3799,SDLEN)),
    to_std_logic_vector(to_signed(5321,SDLEN)),
    to_std_logic_vector(to_signed(6437,SDLEN)),
    to_std_logic_vector(to_signed(7919,SDLEN)),
    to_std_logic_vector(to_signed(11643,SDLEN)),
    to_std_logic_vector(to_signed(15810,SDLEN)),
    to_std_logic_vector(to_signed(16846,SDLEN)),
    to_std_logic_vector(to_signed(18119,SDLEN)),
    to_std_logic_vector(to_signed(18980,SDLEN)),
    to_std_logic_vector(to_signed(3455,SDLEN)),
    to_std_logic_vector(to_signed(4157,SDLEN)),
    to_std_logic_vector(to_signed(6838,SDLEN)),
    to_std_logic_vector(to_signed(8199,SDLEN)),
    to_std_logic_vector(to_signed(9877,SDLEN)),
    to_std_logic_vector(to_signed(12314,SDLEN)),
    to_std_logic_vector(to_signed(15905,SDLEN)),
    to_std_logic_vector(to_signed(16826,SDLEN)),
    to_std_logic_vector(to_signed(19949,SDLEN)),
    to_std_logic_vector(to_signed(20892,SDLEN)),
    to_std_logic_vector(to_signed(3052,SDLEN)),
    to_std_logic_vector(to_signed(3769,SDLEN)),
    to_std_logic_vector(to_signed(4891,SDLEN)),
    to_std_logic_vector(to_signed(5810,SDLEN)),
    to_std_logic_vector(to_signed(6977,SDLEN)),
    to_std_logic_vector(to_signed(10126,SDLEN)),
    to_std_logic_vector(to_signed(14788,SDLEN)),
    to_std_logic_vector(to_signed(15990,SDLEN)),
    to_std_logic_vector(to_signed(19773,SDLEN)),
    to_std_logic_vector(to_signed(20904,SDLEN)),
    to_std_logic_vector(to_signed(3671,SDLEN)),
    to_std_logic_vector(to_signed(4356,SDLEN)),
    to_std_logic_vector(to_signed(5827,SDLEN)),
    to_std_logic_vector(to_signed(6997,SDLEN)),
    to_std_logic_vector(to_signed(8460,SDLEN)),
    to_std_logic_vector(to_signed(12084,SDLEN)),
    to_std_logic_vector(to_signed(14154,SDLEN)),
    to_std_logic_vector(to_signed(14939,SDLEN)),
    to_std_logic_vector(to_signed(19247,SDLEN)),
    to_std_logic_vector(to_signed(20423,SDLEN)),
    to_std_logic_vector(to_signed(2716,SDLEN)),
    to_std_logic_vector(to_signed(3684,SDLEN)),
    to_std_logic_vector(to_signed(5246,SDLEN)),
    to_std_logic_vector(to_signed(6686,SDLEN)),
    to_std_logic_vector(to_signed(8463,SDLEN)),
    to_std_logic_vector(to_signed(10001,SDLEN)),
    to_std_logic_vector(to_signed(12394,SDLEN)),
    to_std_logic_vector(to_signed(14131,SDLEN)),
    to_std_logic_vector(to_signed(16150,SDLEN)),
    to_std_logic_vector(to_signed(19776,SDLEN)),
    to_std_logic_vector(to_signed(1945,SDLEN)),
    to_std_logic_vector(to_signed(2638,SDLEN)),
    to_std_logic_vector(to_signed(4130,SDLEN)),
    to_std_logic_vector(to_signed(7995,SDLEN)),
    to_std_logic_vector(to_signed(14338,SDLEN)),
    to_std_logic_vector(to_signed(15576,SDLEN)),
    to_std_logic_vector(to_signed(17057,SDLEN)),
    to_std_logic_vector(to_signed(18206,SDLEN)),
    to_std_logic_vector(to_signed(20225,SDLEN)),
    to_std_logic_vector(to_signed(20997,SDLEN)),
    to_std_logic_vector(to_signed(2304,SDLEN)),
    to_std_logic_vector(to_signed(2928,SDLEN)),
    to_std_logic_vector(to_signed(4122,SDLEN)),
    to_std_logic_vector(to_signed(4824,SDLEN)),
    to_std_logic_vector(to_signed(5640,SDLEN)),
    to_std_logic_vector(to_signed(13139,SDLEN)),
    to_std_logic_vector(to_signed(15825,SDLEN)),
    to_std_logic_vector(to_signed(16938,SDLEN)),
    to_std_logic_vector(to_signed(20108,SDLEN)),
    to_std_logic_vector(to_signed(21054,SDLEN)),
    to_std_logic_vector(to_signed(1800,SDLEN)),
    to_std_logic_vector(to_signed(2516,SDLEN)),
    to_std_logic_vector(to_signed(3350,SDLEN)),
    to_std_logic_vector(to_signed(5219,SDLEN)),
    to_std_logic_vector(to_signed(13406,SDLEN)),
    to_std_logic_vector(to_signed(15948,SDLEN)),
    to_std_logic_vector(to_signed(17618,SDLEN)),
    to_std_logic_vector(to_signed(18540,SDLEN)),
    to_std_logic_vector(to_signed(20531,SDLEN)),
    to_std_logic_vector(to_signed(21252,SDLEN)),
    to_std_logic_vector(to_signed(1436,SDLEN)),
    to_std_logic_vector(to_signed(2224,SDLEN)),
    to_std_logic_vector(to_signed(2753,SDLEN)),
    to_std_logic_vector(to_signed(4546,SDLEN)),
    to_std_logic_vector(to_signed(9657,SDLEN)),
    to_std_logic_vector(to_signed(11245,SDLEN)),
    to_std_logic_vector(to_signed(15177,SDLEN)),
    to_std_logic_vector(to_signed(16317,SDLEN)),
    to_std_logic_vector(to_signed(17489,SDLEN)),
    to_std_logic_vector(to_signed(19135,SDLEN)),
    to_std_logic_vector(to_signed(2319,SDLEN)),
    to_std_logic_vector(to_signed(2899,SDLEN)),
    to_std_logic_vector(to_signed(4980,SDLEN)),
    to_std_logic_vector(to_signed(6936,SDLEN)),
    to_std_logic_vector(to_signed(8404,SDLEN)),
    to_std_logic_vector(to_signed(13489,SDLEN)),
    to_std_logic_vector(to_signed(15554,SDLEN)),
    to_std_logic_vector(to_signed(16281,SDLEN)),
    to_std_logic_vector(to_signed(20270,SDLEN)),
    to_std_logic_vector(to_signed(20911,SDLEN)),
    to_std_logic_vector(to_signed(2187,SDLEN)),
    to_std_logic_vector(to_signed(2919,SDLEN)),
    to_std_logic_vector(to_signed(4610,SDLEN)),
    to_std_logic_vector(to_signed(5875,SDLEN)),
    to_std_logic_vector(to_signed(7390,SDLEN)),
    to_std_logic_vector(to_signed(12556,SDLEN)),
    to_std_logic_vector(to_signed(14033,SDLEN)),
    to_std_logic_vector(to_signed(16794,SDLEN)),
    to_std_logic_vector(to_signed(20998,SDLEN)),
    to_std_logic_vector(to_signed(21769,SDLEN)),
    to_std_logic_vector(to_signed(2235,SDLEN)),
    to_std_logic_vector(to_signed(2923,SDLEN)),
    to_std_logic_vector(to_signed(5121,SDLEN)),
    to_std_logic_vector(to_signed(6259,SDLEN)),
    to_std_logic_vector(to_signed(8099,SDLEN)),
    to_std_logic_vector(to_signed(13589,SDLEN)),
    to_std_logic_vector(to_signed(15340,SDLEN)),
    to_std_logic_vector(to_signed(16340,SDLEN)),
    to_std_logic_vector(to_signed(17927,SDLEN)),
    to_std_logic_vector(to_signed(20159,SDLEN)),
    to_std_logic_vector(to_signed(1765,SDLEN)),
    to_std_logic_vector(to_signed(2638,SDLEN)),
    to_std_logic_vector(to_signed(3751,SDLEN)),
    to_std_logic_vector(to_signed(5730,SDLEN)),
    to_std_logic_vector(to_signed(7883,SDLEN)),
    to_std_logic_vector(to_signed(10108,SDLEN)),
    to_std_logic_vector(to_signed(13633,SDLEN)),
    to_std_logic_vector(to_signed(15419,SDLEN)),
    to_std_logic_vector(to_signed(16808,SDLEN)),
    to_std_logic_vector(to_signed(18574,SDLEN)),
    to_std_logic_vector(to_signed(3460,SDLEN)),
    to_std_logic_vector(to_signed(5741,SDLEN)),
    to_std_logic_vector(to_signed(9596,SDLEN)),
    to_std_logic_vector(to_signed(11742,SDLEN)),
    to_std_logic_vector(to_signed(14413,SDLEN)),
    to_std_logic_vector(to_signed(16080,SDLEN)),
    to_std_logic_vector(to_signed(18173,SDLEN)),
    to_std_logic_vector(to_signed(19090,SDLEN)),
    to_std_logic_vector(to_signed(20845,SDLEN)),
    to_std_logic_vector(to_signed(21601,SDLEN)),
    to_std_logic_vector(to_signed(3735,SDLEN)),
    to_std_logic_vector(to_signed(4426,SDLEN)),
    to_std_logic_vector(to_signed(6199,SDLEN)),
    to_std_logic_vector(to_signed(7363,SDLEN)),
    to_std_logic_vector(to_signed(9250,SDLEN)),
    to_std_logic_vector(to_signed(14489,SDLEN)),
    to_std_logic_vector(to_signed(16035,SDLEN)),
    to_std_logic_vector(to_signed(17026,SDLEN)),
    to_std_logic_vector(to_signed(19873,SDLEN)),
    to_std_logic_vector(to_signed(20876,SDLEN)),
    to_std_logic_vector(to_signed(3521,SDLEN)),
    to_std_logic_vector(to_signed(4778,SDLEN)),
    to_std_logic_vector(to_signed(6887,SDLEN)),
    to_std_logic_vector(to_signed(8680,SDLEN)),
    to_std_logic_vector(to_signed(12717,SDLEN)),
    to_std_logic_vector(to_signed(14322,SDLEN)),
    to_std_logic_vector(to_signed(15950,SDLEN)),
    to_std_logic_vector(to_signed(18050,SDLEN)),
    to_std_logic_vector(to_signed(20166,SDLEN)),
    to_std_logic_vector(to_signed(21145,SDLEN)),
    to_std_logic_vector(to_signed(2141,SDLEN)),
    to_std_logic_vector(to_signed(2968,SDLEN)),
    to_std_logic_vector(to_signed(6865,SDLEN)),
    to_std_logic_vector(to_signed(8051,SDLEN)),
    to_std_logic_vector(to_signed(10010,SDLEN)),
    to_std_logic_vector(to_signed(13159,SDLEN)),
    to_std_logic_vector(to_signed(14813,SDLEN)),
    to_std_logic_vector(to_signed(15861,SDLEN)),
    to_std_logic_vector(to_signed(17528,SDLEN)),
    to_std_logic_vector(to_signed(18655,SDLEN)),
    to_std_logic_vector(to_signed(4148,SDLEN)),
    to_std_logic_vector(to_signed(6128,SDLEN)),
    to_std_logic_vector(to_signed(9028,SDLEN)),
    to_std_logic_vector(to_signed(10871,SDLEN)),
    to_std_logic_vector(to_signed(12686,SDLEN)),
    to_std_logic_vector(to_signed(14005,SDLEN)),
    to_std_logic_vector(to_signed(15976,SDLEN)),
    to_std_logic_vector(to_signed(17208,SDLEN)),
    to_std_logic_vector(to_signed(19587,SDLEN)),
    to_std_logic_vector(to_signed(20595,SDLEN)),
    to_std_logic_vector(to_signed(4403,SDLEN)),
    to_std_logic_vector(to_signed(5367,SDLEN)),
    to_std_logic_vector(to_signed(6634,SDLEN)),
    to_std_logic_vector(to_signed(8371,SDLEN)),
    to_std_logic_vector(to_signed(10163,SDLEN)),
    to_std_logic_vector(to_signed(11599,SDLEN)),
    to_std_logic_vector(to_signed(14963,SDLEN)),
    to_std_logic_vector(to_signed(16331,SDLEN)),
    to_std_logic_vector(to_signed(17982,SDLEN)),
    to_std_logic_vector(to_signed(18768,SDLEN)),
    to_std_logic_vector(to_signed(4091,SDLEN)),
    to_std_logic_vector(to_signed(5386,SDLEN)),
    to_std_logic_vector(to_signed(6852,SDLEN)),
    to_std_logic_vector(to_signed(8770,SDLEN)),
    to_std_logic_vector(to_signed(11563,SDLEN)),
    to_std_logic_vector(to_signed(13290,SDLEN)),
    to_std_logic_vector(to_signed(15728,SDLEN)),
    to_std_logic_vector(to_signed(16930,SDLEN)),
    to_std_logic_vector(to_signed(19056,SDLEN)),
    to_std_logic_vector(to_signed(20102,SDLEN)),
    to_std_logic_vector(to_signed(2746,SDLEN)),
    to_std_logic_vector(to_signed(3625,SDLEN)),
    to_std_logic_vector(to_signed(5299,SDLEN)),
    to_std_logic_vector(to_signed(7504,SDLEN)),
    to_std_logic_vector(to_signed(10262,SDLEN)),
    to_std_logic_vector(to_signed(11432,SDLEN)),
    to_std_logic_vector(to_signed(13172,SDLEN)),
    to_std_logic_vector(to_signed(15490,SDLEN)),
    to_std_logic_vector(to_signed(16875,SDLEN)),
    to_std_logic_vector(to_signed(17514,SDLEN)),
    to_std_logic_vector(to_signed(2248,SDLEN)),
    to_std_logic_vector(to_signed(3556,SDLEN)),
    to_std_logic_vector(to_signed(8539,SDLEN)),
    to_std_logic_vector(to_signed(10590,SDLEN)),
    to_std_logic_vector(to_signed(12665,SDLEN)),
    to_std_logic_vector(to_signed(14696,SDLEN)),
    to_std_logic_vector(to_signed(16515,SDLEN)),
    to_std_logic_vector(to_signed(17824,SDLEN)),
    to_std_logic_vector(to_signed(20268,SDLEN)),
    to_std_logic_vector(to_signed(21247,SDLEN)),
    to_std_logic_vector(to_signed(1279,SDLEN)),
    to_std_logic_vector(to_signed(1960,SDLEN)),
    to_std_logic_vector(to_signed(3920,SDLEN)),
    to_std_logic_vector(to_signed(7793,SDLEN)),
    to_std_logic_vector(to_signed(10153,SDLEN)),
    to_std_logic_vector(to_signed(14753,SDLEN)),
    to_std_logic_vector(to_signed(16646,SDLEN)),
    to_std_logic_vector(to_signed(18139,SDLEN)),
    to_std_logic_vector(to_signed(20679,SDLEN)),
    to_std_logic_vector(to_signed(21466,SDLEN)),
    to_std_logic_vector(to_signed(2440,SDLEN)),
    to_std_logic_vector(to_signed(3475,SDLEN)),
    to_std_logic_vector(to_signed(6737,SDLEN)),
    to_std_logic_vector(to_signed(8654,SDLEN)),
    to_std_logic_vector(to_signed(12190,SDLEN)),
    to_std_logic_vector(to_signed(14588,SDLEN)),
    to_std_logic_vector(to_signed(17119,SDLEN)),
    to_std_logic_vector(to_signed(17925,SDLEN)),
    to_std_logic_vector(to_signed(19110,SDLEN)),
    to_std_logic_vector(to_signed(19979,SDLEN)),
    to_std_logic_vector(to_signed(1879,SDLEN)),
    to_std_logic_vector(to_signed(2514,SDLEN)),
    to_std_logic_vector(to_signed(4497,SDLEN)),
    to_std_logic_vector(to_signed(7572,SDLEN)),
    to_std_logic_vector(to_signed(10017,SDLEN)),
    to_std_logic_vector(to_signed(14948,SDLEN)),
    to_std_logic_vector(to_signed(16141,SDLEN)),
    to_std_logic_vector(to_signed(16897,SDLEN)),
    to_std_logic_vector(to_signed(18397,SDLEN)),
    to_std_logic_vector(to_signed(19376,SDLEN)),
    to_std_logic_vector(to_signed(2804,SDLEN)),
    to_std_logic_vector(to_signed(3688,SDLEN)),
    to_std_logic_vector(to_signed(7490,SDLEN)),
    to_std_logic_vector(to_signed(10086,SDLEN)),
    to_std_logic_vector(to_signed(11218,SDLEN)),
    to_std_logic_vector(to_signed(12711,SDLEN)),
    to_std_logic_vector(to_signed(16307,SDLEN)),
    to_std_logic_vector(to_signed(17470,SDLEN)),
    to_std_logic_vector(to_signed(20077,SDLEN)),
    to_std_logic_vector(to_signed(21126,SDLEN)),
    to_std_logic_vector(to_signed(2023,SDLEN)),
    to_std_logic_vector(to_signed(2682,SDLEN)),
    to_std_logic_vector(to_signed(3873,SDLEN)),
    to_std_logic_vector(to_signed(8268,SDLEN)),
    to_std_logic_vector(to_signed(10255,SDLEN)),
    to_std_logic_vector(to_signed(11645,SDLEN)),
    to_std_logic_vector(to_signed(15187,SDLEN)),
    to_std_logic_vector(to_signed(17102,SDLEN)),
    to_std_logic_vector(to_signed(18965,SDLEN)),
    to_std_logic_vector(to_signed(19788,SDLEN)),
    to_std_logic_vector(to_signed(2823,SDLEN)),
    to_std_logic_vector(to_signed(3605,SDLEN)),
    to_std_logic_vector(to_signed(5815,SDLEN)),
    to_std_logic_vector(to_signed(8595,SDLEN)),
    to_std_logic_vector(to_signed(10085,SDLEN)),
    to_std_logic_vector(to_signed(11469,SDLEN)),
    to_std_logic_vector(to_signed(16568,SDLEN)),
    to_std_logic_vector(to_signed(17462,SDLEN)),
    to_std_logic_vector(to_signed(18754,SDLEN)),
    to_std_logic_vector(to_signed(19876,SDLEN)),
    to_std_logic_vector(to_signed(2851,SDLEN)),
    to_std_logic_vector(to_signed(3681,SDLEN)),
    to_std_logic_vector(to_signed(5280,SDLEN)),
    to_std_logic_vector(to_signed(7648,SDLEN)),
    to_std_logic_vector(to_signed(9173,SDLEN)),
    to_std_logic_vector(to_signed(10338,SDLEN)),
    to_std_logic_vector(to_signed(14961,SDLEN)),
    to_std_logic_vector(to_signed(16148,SDLEN)),
    to_std_logic_vector(to_signed(17559,SDLEN)),
    to_std_logic_vector(to_signed(18474,SDLEN)),
    to_std_logic_vector(to_signed(1348,SDLEN)),
    to_std_logic_vector(to_signed(2645,SDLEN)),
    to_std_logic_vector(to_signed(5826,SDLEN)),
    to_std_logic_vector(to_signed(8785,SDLEN)),
    to_std_logic_vector(to_signed(10620,SDLEN)),
    to_std_logic_vector(to_signed(12831,SDLEN)),
    to_std_logic_vector(to_signed(16255,SDLEN)),
    to_std_logic_vector(to_signed(18319,SDLEN)),
    to_std_logic_vector(to_signed(21133,SDLEN)),
    to_std_logic_vector(to_signed(22586,SDLEN)),
    to_std_logic_vector(to_signed(2141,SDLEN)),
    to_std_logic_vector(to_signed(3036,SDLEN)),
    to_std_logic_vector(to_signed(4293,SDLEN)),
    to_std_logic_vector(to_signed(6082,SDLEN)),
    to_std_logic_vector(to_signed(7593,SDLEN)),
    to_std_logic_vector(to_signed(10629,SDLEN)),
    to_std_logic_vector(to_signed(17158,SDLEN)),
    to_std_logic_vector(to_signed(18033,SDLEN)),
    to_std_logic_vector(to_signed(21466,SDLEN)),
    to_std_logic_vector(to_signed(22084,SDLEN)),
    to_std_logic_vector(to_signed(1608,SDLEN)),
    to_std_logic_vector(to_signed(2375,SDLEN)),
    to_std_logic_vector(to_signed(3384,SDLEN)),
    to_std_logic_vector(to_signed(6878,SDLEN)),
    to_std_logic_vector(to_signed(9970,SDLEN)),
    to_std_logic_vector(to_signed(11227,SDLEN)),
    to_std_logic_vector(to_signed(16928,SDLEN)),
    to_std_logic_vector(to_signed(17650,SDLEN)),
    to_std_logic_vector(to_signed(20185,SDLEN)),
    to_std_logic_vector(to_signed(21120,SDLEN)),
    to_std_logic_vector(to_signed(2774,SDLEN)),
    to_std_logic_vector(to_signed(3616,SDLEN)),
    to_std_logic_vector(to_signed(5014,SDLEN)),
    to_std_logic_vector(to_signed(6557,SDLEN)),
    to_std_logic_vector(to_signed(7788,SDLEN)),
    to_std_logic_vector(to_signed(8959,SDLEN)),
    to_std_logic_vector(to_signed(17068,SDLEN)),
    to_std_logic_vector(to_signed(18302,SDLEN)),
    to_std_logic_vector(to_signed(19537,SDLEN)),
    to_std_logic_vector(to_signed(20542,SDLEN)),
    to_std_logic_vector(to_signed(1934,SDLEN)),
    to_std_logic_vector(to_signed(4813,SDLEN)),
    to_std_logic_vector(to_signed(6204,SDLEN)),
    to_std_logic_vector(to_signed(7212,SDLEN)),
    to_std_logic_vector(to_signed(8979,SDLEN)),
    to_std_logic_vector(to_signed(11665,SDLEN)),
    to_std_logic_vector(to_signed(15989,SDLEN)),
    to_std_logic_vector(to_signed(17811,SDLEN)),
    to_std_logic_vector(to_signed(20426,SDLEN)),
    to_std_logic_vector(to_signed(21703,SDLEN)),
    to_std_logic_vector(to_signed(2288,SDLEN)),
    to_std_logic_vector(to_signed(3507,SDLEN)),
    to_std_logic_vector(to_signed(5037,SDLEN)),
    to_std_logic_vector(to_signed(6841,SDLEN)),
    to_std_logic_vector(to_signed(8278,SDLEN)),
    to_std_logic_vector(to_signed(9638,SDLEN)),
    to_std_logic_vector(to_signed(15066,SDLEN)),
    to_std_logic_vector(to_signed(16481,SDLEN)),
    to_std_logic_vector(to_signed(21653,SDLEN)),
    to_std_logic_vector(to_signed(22214,SDLEN)),
    to_std_logic_vector(to_signed(2951,SDLEN)),
    to_std_logic_vector(to_signed(3771,SDLEN)),
    to_std_logic_vector(to_signed(4878,SDLEN)),
    to_std_logic_vector(to_signed(7578,SDLEN)),
    to_std_logic_vector(to_signed(9016,SDLEN)),
    to_std_logic_vector(to_signed(10298,SDLEN)),
    to_std_logic_vector(to_signed(14490,SDLEN)),
    to_std_logic_vector(to_signed(15242,SDLEN)),
    to_std_logic_vector(to_signed(20223,SDLEN)),
    to_std_logic_vector(to_signed(20990,SDLEN)),
    to_std_logic_vector(to_signed(3256,SDLEN)),
    to_std_logic_vector(to_signed(4791,SDLEN)),
    to_std_logic_vector(to_signed(6601,SDLEN)),
    to_std_logic_vector(to_signed(7521,SDLEN)),
    to_std_logic_vector(to_signed(8644,SDLEN)),
    to_std_logic_vector(to_signed(9707,SDLEN)),
    to_std_logic_vector(to_signed(13398,SDLEN)),
    to_std_logic_vector(to_signed(16078,SDLEN)),
    to_std_logic_vector(to_signed(19102,SDLEN)),
    to_std_logic_vector(to_signed(20249,SDLEN)),
    to_std_logic_vector(to_signed(1827,SDLEN)),
    to_std_logic_vector(to_signed(2614,SDLEN)),
    to_std_logic_vector(to_signed(3486,SDLEN)),
    to_std_logic_vector(to_signed(6039,SDLEN)),
    to_std_logic_vector(to_signed(12149,SDLEN)),
    to_std_logic_vector(to_signed(13823,SDLEN)),
    to_std_logic_vector(to_signed(16191,SDLEN)),
    to_std_logic_vector(to_signed(17282,SDLEN)),
    to_std_logic_vector(to_signed(21423,SDLEN)),
    to_std_logic_vector(to_signed(22041,SDLEN)),
    to_std_logic_vector(to_signed(1000,SDLEN)),
    to_std_logic_vector(to_signed(1704,SDLEN)),
    to_std_logic_vector(to_signed(3002,SDLEN)),
    to_std_logic_vector(to_signed(6335,SDLEN)),
    to_std_logic_vector(to_signed(8471,SDLEN)),
    to_std_logic_vector(to_signed(10500,SDLEN)),
    to_std_logic_vector(to_signed(14878,SDLEN)),
    to_std_logic_vector(to_signed(16979,SDLEN)),
    to_std_logic_vector(to_signed(20026,SDLEN)),
    to_std_logic_vector(to_signed(22427,SDLEN)),
    to_std_logic_vector(to_signed(1646,SDLEN)),
    to_std_logic_vector(to_signed(2286,SDLEN)),
    to_std_logic_vector(to_signed(3109,SDLEN)),
    to_std_logic_vector(to_signed(7245,SDLEN)),
    to_std_logic_vector(to_signed(11493,SDLEN)),
    to_std_logic_vector(to_signed(12791,SDLEN)),
    to_std_logic_vector(to_signed(16824,SDLEN)),
    to_std_logic_vector(to_signed(17667,SDLEN)),
    to_std_logic_vector(to_signed(18981,SDLEN)),
    to_std_logic_vector(to_signed(20222,SDLEN)),
    to_std_logic_vector(to_signed(1708,SDLEN)),
    to_std_logic_vector(to_signed(2501,SDLEN)),
    to_std_logic_vector(to_signed(3315,SDLEN)),
    to_std_logic_vector(to_signed(6737,SDLEN)),
    to_std_logic_vector(to_signed(8729,SDLEN)),
    to_std_logic_vector(to_signed(9924,SDLEN)),
    to_std_logic_vector(to_signed(16089,SDLEN)),
    to_std_logic_vector(to_signed(17097,SDLEN)),
    to_std_logic_vector(to_signed(18374,SDLEN)),
    to_std_logic_vector(to_signed(19917,SDLEN)),
    to_std_logic_vector(to_signed(2623,SDLEN)),
    to_std_logic_vector(to_signed(3510,SDLEN)),
    to_std_logic_vector(to_signed(4478,SDLEN)),
    to_std_logic_vector(to_signed(5645,SDLEN)),
    to_std_logic_vector(to_signed(9862,SDLEN)),
    to_std_logic_vector(to_signed(11115,SDLEN)),
    to_std_logic_vector(to_signed(15219,SDLEN)),
    to_std_logic_vector(to_signed(18067,SDLEN)),
    to_std_logic_vector(to_signed(19583,SDLEN)),
    to_std_logic_vector(to_signed(20382,SDLEN)),
    to_std_logic_vector(to_signed(2518,SDLEN)),
    to_std_logic_vector(to_signed(3434,SDLEN)),
    to_std_logic_vector(to_signed(4728,SDLEN)),
    to_std_logic_vector(to_signed(6388,SDLEN)),
    to_std_logic_vector(to_signed(8082,SDLEN)),
    to_std_logic_vector(to_signed(9285,SDLEN)),
    to_std_logic_vector(to_signed(13162,SDLEN)),
    to_std_logic_vector(to_signed(18383,SDLEN)),
    to_std_logic_vector(to_signed(19819,SDLEN)),
    to_std_logic_vector(to_signed(20552,SDLEN)),
    to_std_logic_vector(to_signed(1726,SDLEN)),
    to_std_logic_vector(to_signed(2383,SDLEN)),
    to_std_logic_vector(to_signed(4090,SDLEN)),
    to_std_logic_vector(to_signed(6303,SDLEN)),
    to_std_logic_vector(to_signed(7805,SDLEN)),
    to_std_logic_vector(to_signed(12845,SDLEN)),
    to_std_logic_vector(to_signed(14612,SDLEN)),
    to_std_logic_vector(to_signed(17608,SDLEN)),
    to_std_logic_vector(to_signed(19269,SDLEN)),
    to_std_logic_vector(to_signed(20181,SDLEN)),
    to_std_logic_vector(to_signed(2860,SDLEN)),
    to_std_logic_vector(to_signed(3735,SDLEN)),
    to_std_logic_vector(to_signed(4838,SDLEN)),
    to_std_logic_vector(to_signed(6044,SDLEN)),
    to_std_logic_vector(to_signed(7254,SDLEN)),
    to_std_logic_vector(to_signed(8402,SDLEN)),
    to_std_logic_vector(to_signed(14031,SDLEN)),
    to_std_logic_vector(to_signed(16381,SDLEN)),
    to_std_logic_vector(to_signed(18037,SDLEN)),
    to_std_logic_vector(to_signed(19410,SDLEN)),
    to_std_logic_vector(to_signed(4247,SDLEN)),
    to_std_logic_vector(to_signed(5993,SDLEN)),
    to_std_logic_vector(to_signed(7952,SDLEN)),
    to_std_logic_vector(to_signed(9792,SDLEN)),
    to_std_logic_vector(to_signed(12342,SDLEN)),
    to_std_logic_vector(to_signed(14653,SDLEN)),
    to_std_logic_vector(to_signed(17527,SDLEN)),
    to_std_logic_vector(to_signed(18774,SDLEN)),
    to_std_logic_vector(to_signed(20831,SDLEN)),
    to_std_logic_vector(to_signed(21699,SDLEN)),
    to_std_logic_vector(to_signed(3502,SDLEN)),
    to_std_logic_vector(to_signed(4051,SDLEN)),
    to_std_logic_vector(to_signed(5680,SDLEN)),
    to_std_logic_vector(to_signed(6805,SDLEN)),
    to_std_logic_vector(to_signed(8146,SDLEN)),
    to_std_logic_vector(to_signed(11945,SDLEN)),
    to_std_logic_vector(to_signed(16649,SDLEN)),
    to_std_logic_vector(to_signed(17444,SDLEN)),
    to_std_logic_vector(to_signed(20390,SDLEN)),
    to_std_logic_vector(to_signed(21564,SDLEN)),
    to_std_logic_vector(to_signed(3151,SDLEN)),
    to_std_logic_vector(to_signed(4893,SDLEN)),
    to_std_logic_vector(to_signed(5899,SDLEN)),
    to_std_logic_vector(to_signed(7198,SDLEN)),
    to_std_logic_vector(to_signed(11418,SDLEN)),
    to_std_logic_vector(to_signed(13073,SDLEN)),
    to_std_logic_vector(to_signed(15124,SDLEN)),
    to_std_logic_vector(to_signed(17673,SDLEN)),
    to_std_logic_vector(to_signed(20520,SDLEN)),
    to_std_logic_vector(to_signed(21861,SDLEN)),
    to_std_logic_vector(to_signed(3960,SDLEN)),
    to_std_logic_vector(to_signed(4848,SDLEN)),
    to_std_logic_vector(to_signed(5926,SDLEN)),
    to_std_logic_vector(to_signed(7259,SDLEN)),
    to_std_logic_vector(to_signed(8811,SDLEN)),
    to_std_logic_vector(to_signed(10529,SDLEN)),
    to_std_logic_vector(to_signed(15661,SDLEN)),
    to_std_logic_vector(to_signed(16560,SDLEN)),
    to_std_logic_vector(to_signed(18196,SDLEN)),
    to_std_logic_vector(to_signed(20183,SDLEN)),
    to_std_logic_vector(to_signed(4499,SDLEN)),
    to_std_logic_vector(to_signed(6604,SDLEN)),
    to_std_logic_vector(to_signed(8036,SDLEN)),
    to_std_logic_vector(to_signed(9251,SDLEN)),
    to_std_logic_vector(to_signed(10804,SDLEN)),
    to_std_logic_vector(to_signed(12627,SDLEN)),
    to_std_logic_vector(to_signed(15880,SDLEN)),
    to_std_logic_vector(to_signed(17512,SDLEN)),
    to_std_logic_vector(to_signed(20020,SDLEN)),
    to_std_logic_vector(to_signed(21046,SDLEN)),
    to_std_logic_vector(to_signed(4251,SDLEN)),
    to_std_logic_vector(to_signed(5541,SDLEN)),
    to_std_logic_vector(to_signed(6654,SDLEN)),
    to_std_logic_vector(to_signed(8318,SDLEN)),
    to_std_logic_vector(to_signed(9900,SDLEN)),
    to_std_logic_vector(to_signed(11686,SDLEN)),
    to_std_logic_vector(to_signed(15100,SDLEN)),
    to_std_logic_vector(to_signed(17093,SDLEN)),
    to_std_logic_vector(to_signed(20572,SDLEN)),
    to_std_logic_vector(to_signed(21687,SDLEN)),
    to_std_logic_vector(to_signed(3769,SDLEN)),
    to_std_logic_vector(to_signed(5327,SDLEN)),
    to_std_logic_vector(to_signed(7865,SDLEN)),
    to_std_logic_vector(to_signed(9360,SDLEN)),
    to_std_logic_vector(to_signed(10684,SDLEN)),
    to_std_logic_vector(to_signed(11818,SDLEN)),
    to_std_logic_vector(to_signed(13660,SDLEN)),
    to_std_logic_vector(to_signed(15366,SDLEN)),
    to_std_logic_vector(to_signed(18733,SDLEN)),
    to_std_logic_vector(to_signed(19882,SDLEN)),
    to_std_logic_vector(to_signed(3083,SDLEN)),
    to_std_logic_vector(to_signed(3969,SDLEN)),
    to_std_logic_vector(to_signed(6248,SDLEN)),
    to_std_logic_vector(to_signed(8121,SDLEN)),
    to_std_logic_vector(to_signed(9798,SDLEN)),
    to_std_logic_vector(to_signed(10994,SDLEN)),
    to_std_logic_vector(to_signed(12393,SDLEN)),
    to_std_logic_vector(to_signed(13686,SDLEN)),
    to_std_logic_vector(to_signed(17888,SDLEN)),
    to_std_logic_vector(to_signed(19105,SDLEN)),
    to_std_logic_vector(to_signed(2731,SDLEN)),
    to_std_logic_vector(to_signed(4670,SDLEN)),
    to_std_logic_vector(to_signed(7063,SDLEN)),
    to_std_logic_vector(to_signed(9201,SDLEN)),
    to_std_logic_vector(to_signed(11346,SDLEN)),
    to_std_logic_vector(to_signed(13735,SDLEN)),
    to_std_logic_vector(to_signed(16875,SDLEN)),
    to_std_logic_vector(to_signed(18797,SDLEN)),
    to_std_logic_vector(to_signed(20787,SDLEN)),
    to_std_logic_vector(to_signed(22360,SDLEN)),
    to_std_logic_vector(to_signed(1187,SDLEN)),
    to_std_logic_vector(to_signed(2227,SDLEN)),
    to_std_logic_vector(to_signed(4737,SDLEN)),
    to_std_logic_vector(to_signed(7214,SDLEN)),
    to_std_logic_vector(to_signed(9622,SDLEN)),
    to_std_logic_vector(to_signed(12633,SDLEN)),
    to_std_logic_vector(to_signed(15404,SDLEN)),
    to_std_logic_vector(to_signed(17968,SDLEN)),
    to_std_logic_vector(to_signed(20262,SDLEN)),
    to_std_logic_vector(to_signed(23533,SDLEN)),
    to_std_logic_vector(to_signed(1911,SDLEN)),
    to_std_logic_vector(to_signed(2477,SDLEN)),
    to_std_logic_vector(to_signed(3915,SDLEN)),
    to_std_logic_vector(to_signed(10098,SDLEN)),
    to_std_logic_vector(to_signed(11616,SDLEN)),
    to_std_logic_vector(to_signed(12955,SDLEN)),
    to_std_logic_vector(to_signed(16223,SDLEN)),
    to_std_logic_vector(to_signed(17138,SDLEN)),
    to_std_logic_vector(to_signed(19270,SDLEN)),
    to_std_logic_vector(to_signed(20729,SDLEN)),
    to_std_logic_vector(to_signed(1764,SDLEN)),
    to_std_logic_vector(to_signed(2519,SDLEN)),
    to_std_logic_vector(to_signed(3887,SDLEN)),
    to_std_logic_vector(to_signed(6944,SDLEN)),
    to_std_logic_vector(to_signed(9150,SDLEN)),
    to_std_logic_vector(to_signed(12590,SDLEN)),
    to_std_logic_vector(to_signed(16258,SDLEN)),
    to_std_logic_vector(to_signed(16984,SDLEN)),
    to_std_logic_vector(to_signed(17924,SDLEN)),
    to_std_logic_vector(to_signed(18435,SDLEN)),
    to_std_logic_vector(to_signed(1400,SDLEN)),
    to_std_logic_vector(to_signed(3674,SDLEN)),
    to_std_logic_vector(to_signed(7131,SDLEN)),
    to_std_logic_vector(to_signed(8718,SDLEN)),
    to_std_logic_vector(to_signed(10688,SDLEN)),
    to_std_logic_vector(to_signed(12508,SDLEN)),
    to_std_logic_vector(to_signed(15708,SDLEN)),
    to_std_logic_vector(to_signed(17711,SDLEN)),
    to_std_logic_vector(to_signed(19720,SDLEN)),
    to_std_logic_vector(to_signed(21068,SDLEN)),
    to_std_logic_vector(to_signed(2322,SDLEN)),
    to_std_logic_vector(to_signed(3073,SDLEN)),
    to_std_logic_vector(to_signed(4287,SDLEN)),
    to_std_logic_vector(to_signed(8108,SDLEN)),
    to_std_logic_vector(to_signed(9407,SDLEN)),
    to_std_logic_vector(to_signed(10628,SDLEN)),
    to_std_logic_vector(to_signed(15862,SDLEN)),
    to_std_logic_vector(to_signed(16693,SDLEN)),
    to_std_logic_vector(to_signed(19714,SDLEN)),
    to_std_logic_vector(to_signed(21474,SDLEN)),
    to_std_logic_vector(to_signed(2630,SDLEN)),
    to_std_logic_vector(to_signed(3339,SDLEN)),
    to_std_logic_vector(to_signed(4758,SDLEN)),
    to_std_logic_vector(to_signed(8360,SDLEN)),
    to_std_logic_vector(to_signed(10274,SDLEN)),
    to_std_logic_vector(to_signed(11333,SDLEN)),
    to_std_logic_vector(to_signed(12880,SDLEN)),
    to_std_logic_vector(to_signed(17374,SDLEN)),
    to_std_logic_vector(to_signed(19221,SDLEN)),
    to_std_logic_vector(to_signed(19936,SDLEN)),
    to_std_logic_vector(to_signed(1721,SDLEN)),
    to_std_logic_vector(to_signed(2577,SDLEN)),
    to_std_logic_vector(to_signed(5553,SDLEN)),
    to_std_logic_vector(to_signed(7195,SDLEN)),
    to_std_logic_vector(to_signed(8651,SDLEN)),
    to_std_logic_vector(to_signed(10686,SDLEN)),
    to_std_logic_vector(to_signed(15069,SDLEN)),
    to_std_logic_vector(to_signed(16953,SDLEN)),
    to_std_logic_vector(to_signed(18703,SDLEN)),
    to_std_logic_vector(to_signed(19929,SDLEN)),
    to_std_logic_vector(to_signed(-435,SDLEN)),
    to_std_logic_vector(to_signed(-815,SDLEN)),
    to_std_logic_vector(to_signed(-742,SDLEN)),
    to_std_logic_vector(to_signed(1033,SDLEN)),
    to_std_logic_vector(to_signed(-518,SDLEN)),
    to_std_logic_vector(to_signed(582,SDLEN)),
    to_std_logic_vector(to_signed(-1201,SDLEN)),
    to_std_logic_vector(to_signed(829,SDLEN)),
    to_std_logic_vector(to_signed(86,SDLEN)),
    to_std_logic_vector(to_signed(385,SDLEN)),
    to_std_logic_vector(to_signed(-833,SDLEN)),
    to_std_logic_vector(to_signed(-891,SDLEN)),
    to_std_logic_vector(to_signed(463,SDLEN)),
    to_std_logic_vector(to_signed(-8,SDLEN)),
    to_std_logic_vector(to_signed(-1251,SDLEN)),
    to_std_logic_vector(to_signed(1450,SDLEN)),
    to_std_logic_vector(to_signed(72,SDLEN)),
    to_std_logic_vector(to_signed(-231,SDLEN)),
    to_std_logic_vector(to_signed(864,SDLEN)),
    to_std_logic_vector(to_signed(661,SDLEN)),
    to_std_logic_vector(to_signed(-1021,SDLEN)),
    to_std_logic_vector(to_signed(231,SDLEN)),
    to_std_logic_vector(to_signed(-306,SDLEN)),
    to_std_logic_vector(to_signed(321,SDLEN)),
    to_std_logic_vector(to_signed(-220,SDLEN)),
    to_std_logic_vector(to_signed(-163,SDLEN)),
    to_std_logic_vector(to_signed(-526,SDLEN)),
    to_std_logic_vector(to_signed(-754,SDLEN)),
    to_std_logic_vector(to_signed(-1633,SDLEN)),
    to_std_logic_vector(to_signed(267,SDLEN)),
    to_std_logic_vector(to_signed(57,SDLEN)),
    to_std_logic_vector(to_signed(-198,SDLEN)),
    to_std_logic_vector(to_signed(-339,SDLEN)),
    to_std_logic_vector(to_signed(-33,SDLEN)),
    to_std_logic_vector(to_signed(-1468,SDLEN)),
    to_std_logic_vector(to_signed(573,SDLEN)),
    to_std_logic_vector(to_signed(796,SDLEN)),
    to_std_logic_vector(to_signed(-169,SDLEN)),
    to_std_logic_vector(to_signed(-631,SDLEN)),
    to_std_logic_vector(to_signed(816,SDLEN)),
    to_std_logic_vector(to_signed(171,SDLEN)),
    to_std_logic_vector(to_signed(-350,SDLEN)),
    to_std_logic_vector(to_signed(294,SDLEN)),
    to_std_logic_vector(to_signed(1660,SDLEN)),
    to_std_logic_vector(to_signed(453,SDLEN)),
    to_std_logic_vector(to_signed(519,SDLEN)),
    to_std_logic_vector(to_signed(291,SDLEN)),
    to_std_logic_vector(to_signed(159,SDLEN)),
    to_std_logic_vector(to_signed(-640,SDLEN)),
    to_std_logic_vector(to_signed(-1296,SDLEN)),
    to_std_logic_vector(to_signed(-701,SDLEN)),
    to_std_logic_vector(to_signed(-842,SDLEN)),
    to_std_logic_vector(to_signed(-58,SDLEN)),
    to_std_logic_vector(to_signed(950,SDLEN)),
    to_std_logic_vector(to_signed(892,SDLEN)),
    to_std_logic_vector(to_signed(1549,SDLEN)),
    to_std_logic_vector(to_signed(715,SDLEN)),
    to_std_logic_vector(to_signed(527,SDLEN)),
    to_std_logic_vector(to_signed(-714,SDLEN)),
    to_std_logic_vector(to_signed(-193,SDLEN)),
    to_std_logic_vector(to_signed(584,SDLEN)),
    to_std_logic_vector(to_signed(31,SDLEN)),
    to_std_logic_vector(to_signed(-289,SDLEN)),
    to_std_logic_vector(to_signed(356,SDLEN)),
    to_std_logic_vector(to_signed(-333,SDLEN)),
    to_std_logic_vector(to_signed(-457,SDLEN)),
    to_std_logic_vector(to_signed(612,SDLEN)),
    to_std_logic_vector(to_signed(-283,SDLEN)),
    to_std_logic_vector(to_signed(-1381,SDLEN)),
    to_std_logic_vector(to_signed(-741,SDLEN)),
    to_std_logic_vector(to_signed(-109,SDLEN)),
    to_std_logic_vector(to_signed(-808,SDLEN)),
    to_std_logic_vector(to_signed(231,SDLEN)),
    to_std_logic_vector(to_signed(77,SDLEN)),
    to_std_logic_vector(to_signed(-87,SDLEN)),
    to_std_logic_vector(to_signed(-344,SDLEN)),
    to_std_logic_vector(to_signed(1341,SDLEN)),
    to_std_logic_vector(to_signed(1087,SDLEN)),
    to_std_logic_vector(to_signed(-654,SDLEN)),
    to_std_logic_vector(to_signed(-569,SDLEN)),
    to_std_logic_vector(to_signed(-859,SDLEN)),
    to_std_logic_vector(to_signed(1236,SDLEN)),
    to_std_logic_vector(to_signed(550,SDLEN)),
    to_std_logic_vector(to_signed(854,SDLEN)),
    to_std_logic_vector(to_signed(714,SDLEN)),
    to_std_logic_vector(to_signed(-543,SDLEN)),
    to_std_logic_vector(to_signed(-1752,SDLEN)),
    to_std_logic_vector(to_signed(-195,SDLEN)),
    to_std_logic_vector(to_signed(-98,SDLEN)),
    to_std_logic_vector(to_signed(-276,SDLEN)),
    to_std_logic_vector(to_signed(-877,SDLEN)),
    to_std_logic_vector(to_signed(-954,SDLEN)),
    to_std_logic_vector(to_signed(-1248,SDLEN)),
    to_std_logic_vector(to_signed(-299,SDLEN)),
    to_std_logic_vector(to_signed(212,SDLEN)),
    to_std_logic_vector(to_signed(-235,SDLEN)),
    to_std_logic_vector(to_signed(-728,SDLEN)),
    to_std_logic_vector(to_signed(949,SDLEN)),
    to_std_logic_vector(to_signed(1517,SDLEN)),
    to_std_logic_vector(to_signed(895,SDLEN)),
    to_std_logic_vector(to_signed(-77,SDLEN)),
    to_std_logic_vector(to_signed(344,SDLEN)),
    to_std_logic_vector(to_signed(-620,SDLEN)),
    to_std_logic_vector(to_signed(763,SDLEN)),
    to_std_logic_vector(to_signed(413,SDLEN)),
    to_std_logic_vector(to_signed(502,SDLEN)),
    to_std_logic_vector(to_signed(-362,SDLEN)),
    to_std_logic_vector(to_signed(-960,SDLEN)),
    to_std_logic_vector(to_signed(-483,SDLEN)),
    to_std_logic_vector(to_signed(1386,SDLEN)),
    to_std_logic_vector(to_signed(-314,SDLEN)),
    to_std_logic_vector(to_signed(-307,SDLEN)),
    to_std_logic_vector(to_signed(-256,SDLEN)),
    to_std_logic_vector(to_signed(-1260,SDLEN)),
    to_std_logic_vector(to_signed(-429,SDLEN)),
    to_std_logic_vector(to_signed(450,SDLEN)),
    to_std_logic_vector(to_signed(-466,SDLEN)),
    to_std_logic_vector(to_signed(-108,SDLEN)),
    to_std_logic_vector(to_signed(1010,SDLEN)),
    to_std_logic_vector(to_signed(2223,SDLEN)),
    to_std_logic_vector(to_signed(711,SDLEN)),
    to_std_logic_vector(to_signed(693,SDLEN)),
    to_std_logic_vector(to_signed(521,SDLEN)),
    to_std_logic_vector(to_signed(650,SDLEN)),
    to_std_logic_vector(to_signed(1305,SDLEN)),
    to_std_logic_vector(to_signed(-28,SDLEN)),
    to_std_logic_vector(to_signed(-378,SDLEN)),
    to_std_logic_vector(to_signed(744,SDLEN)),
    to_std_logic_vector(to_signed(-1005,SDLEN)),
    to_std_logic_vector(to_signed(240,SDLEN)),
    to_std_logic_vector(to_signed(-112,SDLEN)),
    to_std_logic_vector(to_signed(-271,SDLEN)),
    to_std_logic_vector(to_signed(-500,SDLEN)),
    to_std_logic_vector(to_signed(946,SDLEN)),
    to_std_logic_vector(to_signed(1733,SDLEN)),
    to_std_logic_vector(to_signed(271,SDLEN)),
    to_std_logic_vector(to_signed(-15,SDLEN)),
    to_std_logic_vector(to_signed(909,SDLEN)),
    to_std_logic_vector(to_signed(-259,SDLEN)),
    to_std_logic_vector(to_signed(1688,SDLEN)),
    to_std_logic_vector(to_signed(575,SDLEN)),
    to_std_logic_vector(to_signed(-10,SDLEN)),
    to_std_logic_vector(to_signed(-468,SDLEN)),
    to_std_logic_vector(to_signed(-199,SDLEN)),
    to_std_logic_vector(to_signed(1101,SDLEN)),
    to_std_logic_vector(to_signed(-1011,SDLEN)),
    to_std_logic_vector(to_signed(581,SDLEN)),
    to_std_logic_vector(to_signed(-53,SDLEN)),
    to_std_logic_vector(to_signed(-747,SDLEN)),
    to_std_logic_vector(to_signed(878,SDLEN)),
    to_std_logic_vector(to_signed(145,SDLEN)),
    to_std_logic_vector(to_signed(-285,SDLEN)),
    to_std_logic_vector(to_signed(-1280,SDLEN)),
    to_std_logic_vector(to_signed(-398,SDLEN)),
    to_std_logic_vector(to_signed(36,SDLEN)),
    to_std_logic_vector(to_signed(-498,SDLEN)),
    to_std_logic_vector(to_signed(-1377,SDLEN)),
    to_std_logic_vector(to_signed(18,SDLEN)),
    to_std_logic_vector(to_signed(-444,SDLEN)),
    to_std_logic_vector(to_signed(1483,SDLEN)),
    to_std_logic_vector(to_signed(-1133,SDLEN)),
    to_std_logic_vector(to_signed(-835,SDLEN)),
    to_std_logic_vector(to_signed(1350,SDLEN)),
    to_std_logic_vector(to_signed(1284,SDLEN)),
    to_std_logic_vector(to_signed(-95,SDLEN)),
    to_std_logic_vector(to_signed(1015,SDLEN)),
    to_std_logic_vector(to_signed(-222,SDLEN)),
    to_std_logic_vector(to_signed(443,SDLEN)),
    to_std_logic_vector(to_signed(372,SDLEN)),
    to_std_logic_vector(to_signed(-354,SDLEN)),
    to_std_logic_vector(to_signed(-1459,SDLEN)),
    to_std_logic_vector(to_signed(-1237,SDLEN)),
    to_std_logic_vector(to_signed(416,SDLEN)),
    to_std_logic_vector(to_signed(-213,SDLEN)),
    to_std_logic_vector(to_signed(466,SDLEN)),
    to_std_logic_vector(to_signed(669,SDLEN)),
    to_std_logic_vector(to_signed(659,SDLEN)),
    to_std_logic_vector(to_signed(1640,SDLEN)),
    to_std_logic_vector(to_signed(932,SDLEN)),
    to_std_logic_vector(to_signed(534,SDLEN)),
    to_std_logic_vector(to_signed(-15,SDLEN)),
    to_std_logic_vector(to_signed(66,SDLEN)),
    to_std_logic_vector(to_signed(468,SDLEN)),
    to_std_logic_vector(to_signed(1019,SDLEN)),
    to_std_logic_vector(to_signed(-748,SDLEN)),
    to_std_logic_vector(to_signed(1385,SDLEN)),
    to_std_logic_vector(to_signed(-182,SDLEN)),
    to_std_logic_vector(to_signed(-907,SDLEN)),
    to_std_logic_vector(to_signed(-721,SDLEN)),
    to_std_logic_vector(to_signed(-262,SDLEN)),
    to_std_logic_vector(to_signed(-338,SDLEN)),
    to_std_logic_vector(to_signed(148,SDLEN)),
    to_std_logic_vector(to_signed(1445,SDLEN)),
    to_std_logic_vector(to_signed(75,SDLEN)),
    to_std_logic_vector(to_signed(-760,SDLEN)),
    to_std_logic_vector(to_signed(569,SDLEN)),
    to_std_logic_vector(to_signed(1247,SDLEN)),
    to_std_logic_vector(to_signed(337,SDLEN)),
    to_std_logic_vector(to_signed(416,SDLEN)),
    to_std_logic_vector(to_signed(-121,SDLEN)),
    to_std_logic_vector(to_signed(389,SDLEN)),
    to_std_logic_vector(to_signed(239,SDLEN)),
    to_std_logic_vector(to_signed(1568,SDLEN)),
    to_std_logic_vector(to_signed(981,SDLEN)),
    to_std_logic_vector(to_signed(113,SDLEN)),
    to_std_logic_vector(to_signed(369,SDLEN)),
    to_std_logic_vector(to_signed(-1003,SDLEN)),
    to_std_logic_vector(to_signed(-507,SDLEN)),
    to_std_logic_vector(to_signed(-587,SDLEN)),
    to_std_logic_vector(to_signed(-904,SDLEN)),
    to_std_logic_vector(to_signed(-312,SDLEN)),
    to_std_logic_vector(to_signed(-98,SDLEN)),
    to_std_logic_vector(to_signed(949,SDLEN)),
    to_std_logic_vector(to_signed(31,SDLEN)),
    to_std_logic_vector(to_signed(1104,SDLEN)),
    to_std_logic_vector(to_signed(72,SDLEN)),
    to_std_logic_vector(to_signed(-141,SDLEN)),
    to_std_logic_vector(to_signed(1465,SDLEN)),
    to_std_logic_vector(to_signed(63,SDLEN)),
    to_std_logic_vector(to_signed(-785,SDLEN)),
    to_std_logic_vector(to_signed(1127,SDLEN)),
    to_std_logic_vector(to_signed(584,SDLEN)),
    to_std_logic_vector(to_signed(835,SDLEN)),
    to_std_logic_vector(to_signed(277,SDLEN)),
    to_std_logic_vector(to_signed(-1159,SDLEN)),
    to_std_logic_vector(to_signed(208,SDLEN)),
    to_std_logic_vector(to_signed(301,SDLEN)),
    to_std_logic_vector(to_signed(-882,SDLEN)),
    to_std_logic_vector(to_signed(117,SDLEN)),
    to_std_logic_vector(to_signed(-404,SDLEN)),
    to_std_logic_vector(to_signed(539,SDLEN)),
    to_std_logic_vector(to_signed(-114,SDLEN)),
    to_std_logic_vector(to_signed(856,SDLEN)),
    to_std_logic_vector(to_signed(-493,SDLEN)),
    to_std_logic_vector(to_signed(223,SDLEN)),
    to_std_logic_vector(to_signed(-912,SDLEN)),
    to_std_logic_vector(to_signed(623,SDLEN)),
    to_std_logic_vector(to_signed(-76,SDLEN)),
    to_std_logic_vector(to_signed(276,SDLEN)),
    to_std_logic_vector(to_signed(-440,SDLEN)),
    to_std_logic_vector(to_signed(2197,SDLEN)),
    to_std_logic_vector(to_signed(2337,SDLEN)),
    to_std_logic_vector(to_signed(1268,SDLEN)),
    to_std_logic_vector(to_signed(670,SDLEN)),
    to_std_logic_vector(to_signed(304,SDLEN)),
    to_std_logic_vector(to_signed(-267,SDLEN)),
    to_std_logic_vector(to_signed(-525,SDLEN)),
    to_std_logic_vector(to_signed(140,SDLEN)),
    to_std_logic_vector(to_signed(882,SDLEN)),
    to_std_logic_vector(to_signed(-139,SDLEN)),
    to_std_logic_vector(to_signed(-1596,SDLEN)),
    to_std_logic_vector(to_signed(550,SDLEN)),
    to_std_logic_vector(to_signed(801,SDLEN)),
    to_std_logic_vector(to_signed(-456,SDLEN)),
    to_std_logic_vector(to_signed(-56,SDLEN)),
    to_std_logic_vector(to_signed(-697,SDLEN)),
    to_std_logic_vector(to_signed(865,SDLEN)),
    to_std_logic_vector(to_signed(1060,SDLEN)),
    to_std_logic_vector(to_signed(413,SDLEN)),
    to_std_logic_vector(to_signed(446,SDLEN)),
    to_std_logic_vector(to_signed(1154,SDLEN)),
    to_std_logic_vector(to_signed(593,SDLEN)),
    to_std_logic_vector(to_signed(-77,SDLEN)),
    to_std_logic_vector(to_signed(1237,SDLEN)),
    to_std_logic_vector(to_signed(-31,SDLEN)),
    to_std_logic_vector(to_signed(581,SDLEN)),
    to_std_logic_vector(to_signed(-1037,SDLEN)),
    to_std_logic_vector(to_signed(-895,SDLEN)),
    to_std_logic_vector(to_signed(669,SDLEN)),
    to_std_logic_vector(to_signed(297,SDLEN)),
    to_std_logic_vector(to_signed(397,SDLEN)),
    to_std_logic_vector(to_signed(558,SDLEN)),
    to_std_logic_vector(to_signed(203,SDLEN)),
    to_std_logic_vector(to_signed(-797,SDLEN)),
    to_std_logic_vector(to_signed(-919,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(692,SDLEN)),
    to_std_logic_vector(to_signed(-292,SDLEN)),
    to_std_logic_vector(to_signed(1050,SDLEN)),
    to_std_logic_vector(to_signed(782,SDLEN)),
    to_std_logic_vector(to_signed(334,SDLEN)),
    to_std_logic_vector(to_signed(1475,SDLEN)),
    to_std_logic_vector(to_signed(632,SDLEN)),
    to_std_logic_vector(to_signed(-80,SDLEN)),
    to_std_logic_vector(to_signed(48,SDLEN)),
    to_std_logic_vector(to_signed(-1061,SDLEN)),
    to_std_logic_vector(to_signed(-484,SDLEN)),
    to_std_logic_vector(to_signed(362,SDLEN)),
    to_std_logic_vector(to_signed(-597,SDLEN)),
    to_std_logic_vector(to_signed(-852,SDLEN)),
    to_std_logic_vector(to_signed(-545,SDLEN)),
    to_std_logic_vector(to_signed(-330,SDLEN)),
    to_std_logic_vector(to_signed(-429,SDLEN)),
    to_std_logic_vector(to_signed(-680,SDLEN)),
    to_std_logic_vector(to_signed(1133,SDLEN)),
    to_std_logic_vector(to_signed(-1182,SDLEN)),
    to_std_logic_vector(to_signed(-744,SDLEN)),
    to_std_logic_vector(to_signed(1340,SDLEN)),
    to_std_logic_vector(to_signed(262,SDLEN)),
    to_std_logic_vector(to_signed(63,SDLEN)),
    to_std_logic_vector(to_signed(1320,SDLEN)),
    to_std_logic_vector(to_signed(827,SDLEN)),
    to_std_logic_vector(to_signed(-398,SDLEN)),
    to_std_logic_vector(to_signed(-576,SDLEN)),
    to_std_logic_vector(to_signed(341,SDLEN)),
    to_std_logic_vector(to_signed(-774,SDLEN)),
    to_std_logic_vector(to_signed(-483,SDLEN)),
    to_std_logic_vector(to_signed(-1247,SDLEN)),
    to_std_logic_vector(to_signed(-70,SDLEN)),
    to_std_logic_vector(to_signed(98,SDLEN)),
    to_std_logic_vector(to_signed(-163,SDLEN)),
    to_std_logic_vector(to_signed(674,SDLEN)),
    to_std_logic_vector(to_signed(-11,SDLEN)),
    to_std_logic_vector(to_signed(-886,SDLEN)),
    to_std_logic_vector(to_signed(531,SDLEN)),
    to_std_logic_vector(to_signed(-1125,SDLEN)),
    to_std_logic_vector(to_signed(-265,SDLEN)),
    to_std_logic_vector(to_signed(-242,SDLEN)),
    to_std_logic_vector(to_signed(724,SDLEN)),
    to_std_logic_vector(to_signed(934,SDLEN)),
    to_std_logic_vector(to_signed(8421,SDLEN)),
    to_std_logic_vector(to_signed(9109,SDLEN)),
    to_std_logic_vector(to_signed(9175,SDLEN)),
    to_std_logic_vector(to_signed(8965,SDLEN)),
    to_std_logic_vector(to_signed(9034,SDLEN)),
    to_std_logic_vector(to_signed(9057,SDLEN)),
    to_std_logic_vector(to_signed(8765,SDLEN)),
    to_std_logic_vector(to_signed(8775,SDLEN)),
    to_std_logic_vector(to_signed(9106,SDLEN)),
    to_std_logic_vector(to_signed(8673,SDLEN)),
    to_std_logic_vector(to_signed(7018,SDLEN)),
    to_std_logic_vector(to_signed(7189,SDLEN)),
    to_std_logic_vector(to_signed(7638,SDLEN)),
    to_std_logic_vector(to_signed(7307,SDLEN)),
    to_std_logic_vector(to_signed(7444,SDLEN)),
    to_std_logic_vector(to_signed(7379,SDLEN)),
    to_std_logic_vector(to_signed(7038,SDLEN)),
    to_std_logic_vector(to_signed(6956,SDLEN)),
    to_std_logic_vector(to_signed(6930,SDLEN)),
    to_std_logic_vector(to_signed(6868,SDLEN)),
    to_std_logic_vector(to_signed(5472,SDLEN)),
    to_std_logic_vector(to_signed(4990,SDLEN)),
    to_std_logic_vector(to_signed(5134,SDLEN)),
    to_std_logic_vector(to_signed(5177,SDLEN)),
    to_std_logic_vector(to_signed(5246,SDLEN)),
    to_std_logic_vector(to_signed(5141,SDLEN)),
    to_std_logic_vector(to_signed(5206,SDLEN)),
    to_std_logic_vector(to_signed(5095,SDLEN)),
    to_std_logic_vector(to_signed(4830,SDLEN)),
    to_std_logic_vector(to_signed(5147,SDLEN)),
    to_std_logic_vector(to_signed(4056,SDLEN)),
    to_std_logic_vector(to_signed(3031,SDLEN)),
    to_std_logic_vector(to_signed(2614,SDLEN)),
    to_std_logic_vector(to_signed(3024,SDLEN)),
    to_std_logic_vector(to_signed(2916,SDLEN)),
    to_std_logic_vector(to_signed(2713,SDLEN)),
    to_std_logic_vector(to_signed(3309,SDLEN)),
    to_std_logic_vector(to_signed(3237,SDLEN)),
    to_std_logic_vector(to_signed(2857,SDLEN)),
    to_std_logic_vector(to_signed(3473,SDLEN)),
    to_std_logic_vector(to_signed(7733,SDLEN)),
    to_std_logic_vector(to_signed(7880,SDLEN)),
    to_std_logic_vector(to_signed(8188,SDLEN)),
    to_std_logic_vector(to_signed(8175,SDLEN)),
    to_std_logic_vector(to_signed(8247,SDLEN)),
    to_std_logic_vector(to_signed(8490,SDLEN)),
    to_std_logic_vector(to_signed(8637,SDLEN)),
    to_std_logic_vector(to_signed(8601,SDLEN)),
    to_std_logic_vector(to_signed(8359,SDLEN)),
    to_std_logic_vector(to_signed(7569,SDLEN)),
    to_std_logic_vector(to_signed(4210,SDLEN)),
    to_std_logic_vector(to_signed(3031,SDLEN)),
    to_std_logic_vector(to_signed(2552,SDLEN)),
    to_std_logic_vector(to_signed(3473,SDLEN)),
    to_std_logic_vector(to_signed(3876,SDLEN)),
    to_std_logic_vector(to_signed(3853,SDLEN)),
    to_std_logic_vector(to_signed(4184,SDLEN)),
    to_std_logic_vector(to_signed(4154,SDLEN)),
    to_std_logic_vector(to_signed(3909,SDLEN)),
    to_std_logic_vector(to_signed(3968,SDLEN)),
    to_std_logic_vector(to_signed(3214,SDLEN)),
    to_std_logic_vector(to_signed(1930,SDLEN)),
    to_std_logic_vector(to_signed(1313,SDLEN)),
    to_std_logic_vector(to_signed(2143,SDLEN)),
    to_std_logic_vector(to_signed(2493,SDLEN)),
    to_std_logic_vector(to_signed(2385,SDLEN)),
    to_std_logic_vector(to_signed(2755,SDLEN)),
    to_std_logic_vector(to_signed(2706,SDLEN)),
    to_std_logic_vector(to_signed(2542,SDLEN)),
    to_std_logic_vector(to_signed(2919,SDLEN)),
    to_std_logic_vector(to_signed(3024,SDLEN)),
    to_std_logic_vector(to_signed(1592,SDLEN)),
    to_std_logic_vector(to_signed(940,SDLEN)),
    to_std_logic_vector(to_signed(1631,SDLEN)),
    to_std_logic_vector(to_signed(1723,SDLEN)),
    to_std_logic_vector(to_signed(1579,SDLEN)),
    to_std_logic_vector(to_signed(2034,SDLEN)),
    to_std_logic_vector(to_signed(2084,SDLEN)),
    to_std_logic_vector(to_signed(1913,SDLEN)),
    to_std_logic_vector(to_signed(2601,SDLEN)),
    to_std_logic_vector(to_signed(7798,SDLEN)),
    to_std_logic_vector(to_signed(8447,SDLEN)),
    to_std_logic_vector(to_signed(8205,SDLEN)),
    to_std_logic_vector(to_signed(8293,SDLEN)),
    to_std_logic_vector(to_signed(8126,SDLEN)),
    to_std_logic_vector(to_signed(8477,SDLEN)),
    to_std_logic_vector(to_signed(8447,SDLEN)),
    to_std_logic_vector(to_signed(8703,SDLEN)),
    to_std_logic_vector(to_signed(9043,SDLEN)),
    to_std_logic_vector(to_signed(8604,SDLEN)),
    to_std_logic_vector(to_signed(14585,SDLEN)),
    to_std_logic_vector(to_signed(18333,SDLEN)),
    to_std_logic_vector(to_signed(19772,SDLEN)),
    to_std_logic_vector(to_signed(17344,SDLEN)),
    to_std_logic_vector(to_signed(16426,SDLEN)),
    to_std_logic_vector(to_signed(16459,SDLEN)),
    to_std_logic_vector(to_signed(15155,SDLEN)),
    to_std_logic_vector(to_signed(15220,SDLEN)),
    to_std_logic_vector(to_signed(16043,SDLEN)),
    to_std_logic_vector(to_signed(15708,SDLEN)),
    to_std_logic_vector(to_signed(17210,SDLEN)),
    to_std_logic_vector(to_signed(15888,SDLEN)),
    to_std_logic_vector(to_signed(16357,SDLEN)),
    to_std_logic_vector(to_signed(16183,SDLEN)),
    to_std_logic_vector(to_signed(16516,SDLEN)),
    to_std_logic_vector(to_signed(15833,SDLEN)),
    to_std_logic_vector(to_signed(15888,SDLEN)),
    to_std_logic_vector(to_signed(15421,SDLEN)),
    to_std_logic_vector(to_signed(14840,SDLEN)),
    to_std_logic_vector(to_signed(15597,SDLEN)),
    to_std_logic_vector(to_signed(9202,SDLEN)),
    to_std_logic_vector(to_signed(7320,SDLEN)),
    to_std_logic_vector(to_signed(6788,SDLEN)),
    to_std_logic_vector(to_signed(7738,SDLEN)),
    to_std_logic_vector(to_signed(8170,SDLEN)),
    to_std_logic_vector(to_signed(8154,SDLEN)),
    to_std_logic_vector(to_signed(8856,SDLEN)),
    to_std_logic_vector(to_signed(8818,SDLEN)),
    to_std_logic_vector(to_signed(8366,SDLEN)),
    to_std_logic_vector(to_signed(8544,SDLEN)),
    to_std_logic_vector(to_signed(29443,SDLEN)),
    to_std_logic_vector(to_signed(25207,SDLEN)),
    to_std_logic_vector(to_signed(14701,SDLEN)),
    to_std_logic_vector(to_signed(3143,SDLEN)),
    to_std_logic_vector(to_signed(-4402,SDLEN)),
    to_std_logic_vector(to_signed(-5850,SDLEN)),
    to_std_logic_vector(to_signed(-2783,SDLEN)),
    to_std_logic_vector(to_signed(1211,SDLEN)),
    to_std_logic_vector(to_signed(3130,SDLEN)),
    to_std_logic_vector(to_signed(2259,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(-1652,SDLEN)),
    to_std_logic_vector(to_signed(-1666,SDLEN)),
    to_std_logic_vector(to_signed(-464,SDLEN)),
    to_std_logic_vector(to_signed(756,SDLEN)),
    to_std_logic_vector(to_signed(1099,SDLEN)),
    to_std_logic_vector(to_signed(550,SDLEN)),
    to_std_logic_vector(to_signed(-245,SDLEN)),
    to_std_logic_vector(to_signed(-634,SDLEN)),
    to_std_logic_vector(to_signed(-451,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(308,SDLEN)),
    to_std_logic_vector(to_signed(296,SDLEN)),
    to_std_logic_vector(to_signed(78,SDLEN)),
    to_std_logic_vector(to_signed(-120,SDLEN)),
    to_std_logic_vector(to_signed(-165,SDLEN)),
    to_std_logic_vector(to_signed(-79,SDLEN)),
    to_std_logic_vector(to_signed(34,SDLEN)),
    to_std_logic_vector(to_signed(91,SDLEN)),
    to_std_logic_vector(to_signed(70,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(5571,SDLEN)),
    to_std_logic_vector(to_signed(4751,SDLEN)),
    to_std_logic_vector(to_signed(2785,SDLEN)),
    to_std_logic_vector(to_signed(1556,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1516,SDLEN)),
    to_std_logic_vector(to_signed(1551,SDLEN)),
    to_std_logic_vector(to_signed(2425,SDLEN)),
    to_std_logic_vector(to_signed(1831,SDLEN)),
    to_std_logic_vector(to_signed(5022,SDLEN)),
    to_std_logic_vector(to_signed(57,SDLEN)),
    to_std_logic_vector(to_signed(5404,SDLEN)),
    to_std_logic_vector(to_signed(1921,SDLEN)),
    to_std_logic_vector(to_signed(9291,SDLEN)),
    to_std_logic_vector(to_signed(3242,SDLEN)),
    to_std_logic_vector(to_signed(9949,SDLEN)),
    to_std_logic_vector(to_signed(356,SDLEN)),
    to_std_logic_vector(to_signed(14756,SDLEN)),
    to_std_logic_vector(to_signed(2678,SDLEN)),
    to_std_logic_vector(to_signed(27162,SDLEN)),
    to_std_logic_vector(to_signed(826,SDLEN)),
    to_std_logic_vector(to_signed(2005,SDLEN)),
    to_std_logic_vector(to_signed(1994,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(5142,SDLEN)),
    to_std_logic_vector(to_signed(592,SDLEN)),
    to_std_logic_vector(to_signed(6160,SDLEN)),
    to_std_logic_vector(to_signed(2395,SDLEN)),
    to_std_logic_vector(to_signed(8091,SDLEN)),
    to_std_logic_vector(to_signed(4861,SDLEN)),
    to_std_logic_vector(to_signed(9120,SDLEN)),
    to_std_logic_vector(to_signed(525,SDLEN)),
    to_std_logic_vector(to_signed(10573,SDLEN)),
    to_std_logic_vector(to_signed(2966,SDLEN)),
    to_std_logic_vector(to_signed(11569,SDLEN)),
    to_std_logic_vector(to_signed(1196,SDLEN)),
    to_std_logic_vector(to_signed(13260,SDLEN)),
    to_std_logic_vector(to_signed(3256,SDLEN)),
    to_std_logic_vector(to_signed(14194,SDLEN)),
    to_std_logic_vector(to_signed(1630,SDLEN)),
    to_std_logic_vector(to_signed(15132,SDLEN)),
    to_std_logic_vector(to_signed(4914,SDLEN)),
    to_std_logic_vector(to_signed(15161,SDLEN)),
    to_std_logic_vector(to_signed(14276,SDLEN)),
    to_std_logic_vector(to_signed(15434,SDLEN)),
    to_std_logic_vector(to_signed(237,SDLEN)),
    to_std_logic_vector(to_signed(16112,SDLEN)),
    to_std_logic_vector(to_signed(3392,SDLEN)),
    to_std_logic_vector(to_signed(17299,SDLEN)),
    to_std_logic_vector(to_signed(1861,SDLEN)),
    to_std_logic_vector(to_signed(18973,SDLEN)),
    to_std_logic_vector(to_signed(5935,SDLEN)),
    to_std_logic_vector(to_signed(5,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(4,SDLEN)),
    to_std_logic_vector(to_signed(7,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(6,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(4,SDLEN)),
    to_std_logic_vector(to_signed(6,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(12,SDLEN)),
    to_std_logic_vector(to_signed(14,SDLEN)),
    to_std_logic_vector(to_signed(8,SDLEN)),
    to_std_logic_vector(to_signed(10,SDLEN)),
    to_std_logic_vector(to_signed(15,SDLEN)),
    to_std_logic_vector(to_signed(11,SDLEN)),
    to_std_logic_vector(to_signed(9,SDLEN)),
    to_std_logic_vector(to_signed(13,SDLEN)),
    to_std_logic_vector(to_signed(7,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(5,SDLEN)),
    to_std_logic_vector(to_signed(31881,SDLEN)),
    to_std_logic_vector(to_signed(26416,SDLEN)),
    to_std_logic_vector(to_signed(31548,SDLEN)),
    to_std_logic_vector(to_signed(27816,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(10808,SDLEN)),
    to_std_logic_vector(to_signed(12374,SDLEN)),
    to_std_logic_vector(to_signed(19778,SDLEN)),
    to_std_logic_vector(to_signed(32567,SDLEN)),
    to_std_logic_vector(to_signed(14087,SDLEN)),
    to_std_logic_vector(to_signed(16188,SDLEN)),
    to_std_logic_vector(to_signed(20274,SDLEN)),
    to_std_logic_vector(to_signed(21321,SDLEN)),
    to_std_logic_vector(to_signed(23525,SDLEN)),
    to_std_logic_vector(to_signed(25232,SDLEN)),
    to_std_logic_vector(to_signed(27873,SDLEN)),
    to_std_logic_vector(to_signed(30542,SDLEN)),
    to_std_logic_vector(to_signed(5,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(7,SDLEN)),
    to_std_logic_vector(to_signed(4,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(6,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(14,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(13,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(15,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(12,SDLEN)),
    to_std_logic_vector(to_signed(6,SDLEN)),
    to_std_logic_vector(to_signed(10,SDLEN)),
    to_std_logic_vector(to_signed(7,SDLEN)),
    to_std_logic_vector(to_signed(9,SDLEN)),
    to_std_logic_vector(to_signed(4,SDLEN)),
    to_std_logic_vector(to_signed(11,SDLEN)),
    to_std_logic_vector(to_signed(5,SDLEN)),
    to_std_logic_vector(to_signed(8,SDLEN)),
    to_std_logic_vector(to_signed(7699,SDLEN)),
    to_std_logic_vector(to_signed(-15398,SDLEN)),
    to_std_logic_vector(to_signed(7699,SDLEN)),
    to_std_logic_vector(to_signed(8192,SDLEN)),
    to_std_logic_vector(to_signed(15836,SDLEN)),
    to_std_logic_vector(to_signed(-7667,SDLEN)),
    to_std_logic_vector(to_signed(1899,SDLEN)),
    to_std_logic_vector(to_signed(-3798,SDLEN)),
    to_std_logic_vector(to_signed(1899,SDLEN)),
    to_std_logic_vector(to_signed(4096,SDLEN)),
    to_std_logic_vector(to_signed(7807,SDLEN)),
    to_std_logic_vector(to_signed(-3733,SDLEN)),
    to_std_logic_vector(to_signed(8,SDLEN)),
    to_std_logic_vector(to_signed(10,SDLEN)),
    to_std_logic_vector(to_signed(8,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(13,SDLEN)),
    to_std_logic_vector(to_signed(4,SDLEN)),
    to_std_logic_vector(to_signed(7,SDLEN)),
    to_std_logic_vector(to_signed(5,SDLEN)),
    to_std_logic_vector(to_signed(13,SDLEN)),
    to_std_logic_vector(to_signed(4,SDLEN)),
    to_std_logic_vector(to_signed(7,SDLEN)),
    to_std_logic_vector(to_signed(16384,SDLEN)),
    to_std_logic_vector(to_signed(16743,SDLEN)),
    to_std_logic_vector(to_signed(17109,SDLEN)),
    to_std_logic_vector(to_signed(17484,SDLEN)),
    to_std_logic_vector(to_signed(17867,SDLEN)),
    to_std_logic_vector(to_signed(18258,SDLEN)),
    to_std_logic_vector(to_signed(18658,SDLEN)),
    to_std_logic_vector(to_signed(19066,SDLEN)),
    to_std_logic_vector(to_signed(19484,SDLEN)),
    to_std_logic_vector(to_signed(19911,SDLEN)),
    to_std_logic_vector(to_signed(20347,SDLEN)),
    to_std_logic_vector(to_signed(20792,SDLEN)),
    to_std_logic_vector(to_signed(21247,SDLEN)),
    to_std_logic_vector(to_signed(21713,SDLEN)),
    to_std_logic_vector(to_signed(22188,SDLEN)),
    to_std_logic_vector(to_signed(22674,SDLEN)),
    to_std_logic_vector(to_signed(23170,SDLEN)),
    to_std_logic_vector(to_signed(23678,SDLEN)),
    to_std_logic_vector(to_signed(24196,SDLEN)),
    to_std_logic_vector(to_signed(24726,SDLEN)),
    to_std_logic_vector(to_signed(25268,SDLEN)),
    to_std_logic_vector(to_signed(25821,SDLEN)),
    to_std_logic_vector(to_signed(26386,SDLEN)),
    to_std_logic_vector(to_signed(26964,SDLEN)),
    to_std_logic_vector(to_signed(27554,SDLEN)),
    to_std_logic_vector(to_signed(28158,SDLEN)),
    to_std_logic_vector(to_signed(28774,SDLEN)),
    to_std_logic_vector(to_signed(29405,SDLEN)),
    to_std_logic_vector(to_signed(30048,SDLEN)),
    to_std_logic_vector(to_signed(30706,SDLEN)),
    to_std_logic_vector(to_signed(31379,SDLEN)),
    to_std_logic_vector(to_signed(32066,SDLEN)),
    to_std_logic_vector(to_signed(32767,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(1455,SDLEN)),
    to_std_logic_vector(to_signed(2866,SDLEN)),
    to_std_logic_vector(to_signed(4236,SDLEN)),
    to_std_logic_vector(to_signed(5568,SDLEN)),
    to_std_logic_vector(to_signed(6863,SDLEN)),
    to_std_logic_vector(to_signed(8124,SDLEN)),
    to_std_logic_vector(to_signed(9352,SDLEN)),
    to_std_logic_vector(to_signed(10549,SDLEN)),
    to_std_logic_vector(to_signed(11716,SDLEN)),
    to_std_logic_vector(to_signed(12855,SDLEN)),
    to_std_logic_vector(to_signed(13967,SDLEN)),
    to_std_logic_vector(to_signed(15054,SDLEN)),
    to_std_logic_vector(to_signed(16117,SDLEN)),
    to_std_logic_vector(to_signed(17156,SDLEN)),
    to_std_logic_vector(to_signed(18172,SDLEN)),
    to_std_logic_vector(to_signed(19167,SDLEN)),
    to_std_logic_vector(to_signed(20142,SDLEN)),
    to_std_logic_vector(to_signed(21097,SDLEN)),
    to_std_logic_vector(to_signed(22033,SDLEN)),
    to_std_logic_vector(to_signed(22951,SDLEN)),
    to_std_logic_vector(to_signed(23852,SDLEN)),
    to_std_logic_vector(to_signed(24735,SDLEN)),
    to_std_logic_vector(to_signed(25603,SDLEN)),
    to_std_logic_vector(to_signed(26455,SDLEN)),
    to_std_logic_vector(to_signed(27291,SDLEN)),
    to_std_logic_vector(to_signed(28113,SDLEN)),
    to_std_logic_vector(to_signed(28922,SDLEN)),
    to_std_logic_vector(to_signed(29716,SDLEN)),
    to_std_logic_vector(to_signed(30497,SDLEN)),
    to_std_logic_vector(to_signed(31266,SDLEN)),
    to_std_logic_vector(to_signed(32023,SDLEN)),
    to_std_logic_vector(to_signed(32767,SDLEN)),
    to_std_logic_vector(to_signed(32767,SDLEN)),
    to_std_logic_vector(to_signed(31790,SDLEN)),
    to_std_logic_vector(to_signed(30894,SDLEN)),
    to_std_logic_vector(to_signed(30070,SDLEN)),
    to_std_logic_vector(to_signed(29309,SDLEN)),
    to_std_logic_vector(to_signed(28602,SDLEN)),
    to_std_logic_vector(to_signed(27945,SDLEN)),
    to_std_logic_vector(to_signed(27330,SDLEN)),
    to_std_logic_vector(to_signed(26755,SDLEN)),
    to_std_logic_vector(to_signed(26214,SDLEN)),
    to_std_logic_vector(to_signed(25705,SDLEN)),
    to_std_logic_vector(to_signed(25225,SDLEN)),
    to_std_logic_vector(to_signed(24770,SDLEN)),
    to_std_logic_vector(to_signed(24339,SDLEN)),
    to_std_logic_vector(to_signed(23930,SDLEN)),
    to_std_logic_vector(to_signed(23541,SDLEN)),
    to_std_logic_vector(to_signed(23170,SDLEN)),
    to_std_logic_vector(to_signed(22817,SDLEN)),
    to_std_logic_vector(to_signed(22479,SDLEN)),
    to_std_logic_vector(to_signed(22155,SDLEN)),
    to_std_logic_vector(to_signed(21845,SDLEN)),
    to_std_logic_vector(to_signed(21548,SDLEN)),
    to_std_logic_vector(to_signed(21263,SDLEN)),
    to_std_logic_vector(to_signed(20988,SDLEN)),
    to_std_logic_vector(to_signed(20724,SDLEN)),
    to_std_logic_vector(to_signed(20470,SDLEN)),
    to_std_logic_vector(to_signed(20225,SDLEN)),
    to_std_logic_vector(to_signed(19988,SDLEN)),
    to_std_logic_vector(to_signed(19760,SDLEN)),
    to_std_logic_vector(to_signed(19539,SDLEN)),
    to_std_logic_vector(to_signed(19326,SDLEN)),
    to_std_logic_vector(to_signed(19119,SDLEN)),
    to_std_logic_vector(to_signed(18919,SDLEN)),
    to_std_logic_vector(to_signed(18725,SDLEN)),
    to_std_logic_vector(to_signed(18536,SDLEN)),
    to_std_logic_vector(to_signed(18354,SDLEN)),
    to_std_logic_vector(to_signed(18176,SDLEN)),
    to_std_logic_vector(to_signed(18004,SDLEN)),
    to_std_logic_vector(to_signed(17837,SDLEN)),
    to_std_logic_vector(to_signed(17674,SDLEN)),
    to_std_logic_vector(to_signed(17515,SDLEN)),
    to_std_logic_vector(to_signed(17361,SDLEN)),
    to_std_logic_vector(to_signed(17211,SDLEN)),
    to_std_logic_vector(to_signed(17064,SDLEN)),
    to_std_logic_vector(to_signed(16921,SDLEN)),
    to_std_logic_vector(to_signed(16782,SDLEN)),
    to_std_logic_vector(to_signed(16646,SDLEN)),
    to_std_logic_vector(to_signed(16514,SDLEN)),
    to_std_logic_vector(to_signed(16384,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(32760,SDLEN)),
    to_std_logic_vector(to_signed(32703,SDLEN)),
    to_std_logic_vector(to_signed(32509,SDLEN)),
    to_std_logic_vector(to_signed(32187,SDLEN)),
    to_std_logic_vector(to_signed(31738,SDLEN)),
    to_std_logic_vector(to_signed(31164,SDLEN)),
    to_std_logic_vector(to_signed(30466,SDLEN)),
    to_std_logic_vector(to_signed(29649,SDLEN)),
    to_std_logic_vector(to_signed(28714,SDLEN)),
    to_std_logic_vector(to_signed(27666,SDLEN)),
    to_std_logic_vector(to_signed(26509,SDLEN)),
    to_std_logic_vector(to_signed(25248,SDLEN)),
    to_std_logic_vector(to_signed(23886,SDLEN)),
    to_std_logic_vector(to_signed(22431,SDLEN)),
    to_std_logic_vector(to_signed(20887,SDLEN)),
    to_std_logic_vector(to_signed(19260,SDLEN)),
    to_std_logic_vector(to_signed(17557,SDLEN)),
    to_std_logic_vector(to_signed(15786,SDLEN)),
    to_std_logic_vector(to_signed(13951,SDLEN)),
    to_std_logic_vector(to_signed(12062,SDLEN)),
    to_std_logic_vector(to_signed(10125,SDLEN)),
    to_std_logic_vector(to_signed(8149,SDLEN)),
    to_std_logic_vector(to_signed(6140,SDLEN)),
    to_std_logic_vector(to_signed(4106,SDLEN)),
    to_std_logic_vector(to_signed(2057,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(-2057,SDLEN)),
    to_std_logic_vector(to_signed(-4106,SDLEN)),
    to_std_logic_vector(to_signed(-6140,SDLEN)),
    to_std_logic_vector(to_signed(-8149,SDLEN)),
    to_std_logic_vector(to_signed(-10125,SDLEN)),
    to_std_logic_vector(to_signed(-12062,SDLEN)),
    to_std_logic_vector(to_signed(-13951,SDLEN)),
    to_std_logic_vector(to_signed(-15786,SDLEN)),
    to_std_logic_vector(to_signed(-17557,SDLEN)),
    to_std_logic_vector(to_signed(-19260,SDLEN)),
    to_std_logic_vector(to_signed(-20887,SDLEN)),
    to_std_logic_vector(to_signed(-22431,SDLEN)),
    to_std_logic_vector(to_signed(-23886,SDLEN)),
    to_std_logic_vector(to_signed(-25248,SDLEN)),
    to_std_logic_vector(to_signed(-26509,SDLEN)),
    to_std_logic_vector(to_signed(-27666,SDLEN)),
    to_std_logic_vector(to_signed(-28714,SDLEN)),
    to_std_logic_vector(to_signed(-29649,SDLEN)),
    to_std_logic_vector(to_signed(-30466,SDLEN)),
    to_std_logic_vector(to_signed(-31164,SDLEN)),
    to_std_logic_vector(to_signed(-31738,SDLEN)),
    to_std_logic_vector(to_signed(-32187,SDLEN)),
    to_std_logic_vector(to_signed(-32509,SDLEN)),
    to_std_logic_vector(to_signed(-32703,SDLEN)),
    to_std_logic_vector(to_signed(-32760,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN))
  );

--END;

end G729A_ASIP_ROMD_PKG;

package body G729A_ASIP_ROMD_PKG is

end G729A_ASIP_ROMD_PKG;
