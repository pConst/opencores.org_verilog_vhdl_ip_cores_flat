-----------------------------------------------------------------------
----                                                               ----
---- Montgomery modular multiplier and exponentiator               ----
----                                                               ----
---- This file is part of the Montgomery modular multiplier        ----
---- and exponentiator project                                     ----
---- http://opencores.org/project,mod_mult_exp                     ----
----                                                               ----
---- Description:                                                  ----
----   This is TestBench for the Montgomery modular multiplier     ----
----   with the 512 bit width.                                     ----
----   it takes two nubers and modulus as the input and results    ----
----   the Montgomery product A*B*(R^{-1}) mod M                   ----
----   where R^{-1} is the modular multiplicative inverse.         ----
----   R*R^{-1} == 1 mod M                                         ----
----   R = 2^word_length mod M                                     ----
----               and word_length is the binary width of the      ----
----               operated word (in this case 512 bit)            ----
---- To Do:                                                        ----
----                                                               ----
---- Author(s):                                                    ----
---- - Krzysztof Gajewski, gajos@opencores.org                     ----
----                       k.gajewski@gmail.com                    ----
----                                                               ----
-----------------------------------------------------------------------
----                                                               ----
---- Copyright (C) 2014 Authors and OPENCORES.ORG                  ----
----                                                               ----
---- This source file may be used and distributed without          ----
---- restriction provided that this copyright statement is not     ----
---- removed from the file and that any derivative work contains   ----
---- the original copyright notice and the associated disclaimer.  ----
----                                                               ----
---- This source file is free software; you can redistribute it    ----
---- and-or modify it under the terms of the GNU Lesser General    ----
---- Public License as published by the Free Software Foundation;  ----
---- either version 2.1 of the License, or (at your option) any    ----
---- later version.                                                ----
----                                                               ----
---- This source is distributed in the hope that it will be        ----
---- useful, but WITHOUT ANY WARRANTY; without even the implied    ----
---- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR       ----
---- PURPOSE. See the GNU Lesser General Public License for more   ----
---- details.                                                      ----
----                                                               ----
---- You should have received a copy of the GNU Lesser General     ----
---- Public License along with this source; if not, download it    ----
---- from http://www.opencores.org/lgpl.shtml                      ----
----                                                               ----
-----------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY ModularMultiplierIterative512bitTB IS
END ModularMultiplierIterative512bitTB;
 
ARCHITECTURE behavior OF ModularMultiplierIterative512bitTB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT ModularMultiplierIterative
    PORT(
         A       : in  STD_LOGIC_VECTOR(511 downto 0);
         B       : in  STD_LOGIC_VECTOR(511 downto 0);
         M       : in  STD_LOGIC_VECTOR(511 downto 0);
         start   : in  STD_LOGIC;
         product : out STD_LOGIC_VECTOR(511 downto 0);
         ready   : out STD_LOGIC;
         clk     : in  STD_LOGIC
        );
    END COMPONENT;
    

   --Inputs
   signal A     : STD_LOGIC_VECTOR(511 downto 0) := (others => '0');
   signal B     : STD_LOGIC_VECTOR(511 downto 0) := (others => '0');
   signal M     : STD_LOGIC_VECTOR(511 downto 0) := (others => '0');
   signal start : STD_LOGIC := '0';
   signal clk   : STD_LOGIC := '0';

 	--Outputs
   signal product : STD_LOGIC_VECTOR(511 downto 0);
   signal ready   : STD_LOGIC;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: ModularMultiplierIterative PORT MAP (
          A => A,
          B => B,
          M => M,
          start => start,
          product => product,
          ready => ready,
          clk => clk
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      
		start <= '0';
      wait for 100 ns;	

---- Preparation for test case 1 -----------------
--    A = 1135574785903187283000914738069914842639275616893687122668359807022003618585980215260939798952644749528921700342000274265548842002316414917974647561961683 in decimal
--    B = 97927786390663519429528993360368267006249228136794892056090651513080073109454331808866772457049032741774590681339704155886317906072752116837364369820881 in decimal
--    M = 3351951982485649274893506249551461531869841455148098344430890360930446855046914914263767984168972974033957028381338463851007479808527777429670210341401251 in decimal
--    expected_result = 2228133496571818711622350692880669459929128102839647013792122413518929533298354919965858625663488002993791315812426542313874032336596139553001249634708855 in decimal,  
--               in hex 2a8ae3c12ae96d6babce2e342ec7beeff5754a14e7c8e6057eeebf6dc1cb12145e26e97c874f8e05cfa6fcaf83240f90d2fd21b3f41016b74607c143e49eed77
--    mod(
--        1135574785903187283000914738069914842639275616893687122668359807022003618585980215260939798952644749528921700342000274265548842002316414917974647561961683 * 
--        97927786390663519429528993360368267006249228136794892056090651513080073109454331808866772457049032741774590681339704155886317906072752116837364369820881 * 
--        2591367877621154684380773880291249237701602230100736077754314629198930824379666744084279080961590867282481555124997788427853751639203524473059719065731751 , 
--        3351951982485649274893506249551461531869841455148098344430890360930446855046914914263767984168972974033957028381338463851007479808527777429670210341401251 ) = 
--        = 2228133496571818711622350692880669459929128102839647013792122413518929533298354919965858625663488002993791315812426542313874032336596139553001249634708855
--    where 2591367877621154684380773880291249237701602230100736077754314629198930824379666744084279080961590867282481555124997788427853751639203524473059719065731751 is the inverse modulus
--------------------------------------------------
      
      start <= '1';
      --    A = 1135574785903187283000914738069914842639275616893687122668359807022003618585980215260939798952644749528921700342000274265548842002316414917974647561961683 in decimal
      A <=  "00010101101011101001001011101101001001011100110110111011001010010100010110000100000101001010110100011010001010001111101000110101111101011011111111000011000100011101011111100001111011111110110110111010011101010011111001001000110011001110111000011110100111111111000111010001011000000111000101000100010010011011111101101111100001011010000011100011111111100000011110000100010101001000101100111100010001100001101011000101111110111111001010001011011110100001110000111100100000111111010011011111111101101100000011010011";
      --    B = 97927786390663519429528993360368267006249228136794892056090651513080073109454331808866772457049032741774590681339704155886317906072752116837364369820881 in decimal
	  B <=  "00000001110111101010100100111010100000100100111111101001100100111011001111000010101011111001001001110011011010010100101000100010110011011101111000010011100100101000011010000110110010101101101100000111101000001111010101000110100001100011101110100011100111101100000001000110010110111001110111111110101000001110001000011001000001000000111100000001100110000100011100010011101110010100111110010111110001000110111010010010101101001111110000111001110000100111111111100011011101100000011110100100100000011000110011010001";
      --    M = 3351951982485649274893506249551461531869841455148098344430890360930446855046914914263767984168972974033957028381338463851007479808527777429670210341401251 in decimal
      M <=  "01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001010010010100100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110101111001111111011110110110111001010100011";
	  
	  --wait for 600*clk_period;
      --    Result = 2228133496571818711622350692880669459929128102839647013792122413518929533298354919965858625663488002993791315812426542313874032336596139553001249634708855 in decimal		
	  
	  wait until ready = '1' and clk = '0';
		
	  if product /= x"2a8ae3c12ae96d6babce2e342ec7beeff5754a14e7c8e6057eeebf6dc1cb12145e26e97c874f8e05cfa6fcaf83240f90d2fd21b3f41016b74607c143e49eed77" then
        report "RESULT MISMATCH! Test case 1 failed" severity ERROR;
		assert false severity failure;
	  else
		report "Test case 1 successful" severity note;	
	  end if; 
	  
	  start <= '0';

---- Preparation for test case 2 -----------------
--    A = 3351951982485649274893506249551461531869841455148098344430890360930441007518386744200468574541725856922507964546621512713438470702986642486608412251521039 in decimal
--    B = 97927786390663519429528993360368267006249228136794892056090651513080073109454331808866772457049032741774590681339704155886317906072752116837364369820881 in decimal
--    M = 6703903964971298549787012499102923063739682910296196688861780721860882015036773488400937149083451713845015929093243025426876941405973284973216824503042159 in decimal
--    expected_result = 5770539552593938046267215339235143056108840937616962443047031076129629580294766891795665005337423591502330655021878623252853392851503861478061794255888635 in decimal,  
--               in hex 6e2dcf4e2226cb7a14afa007b0bafdf50d573776681c0cca8d7ff56515076baffd05eaa8ee73d63874a1df6d13e2bbc0aeb6dcd21d8ee10613df1e2e5e02e0fb
--    mod(
--        3351951982485649274893506249551461531869841455148098344430890360930441007518386744200468574541725856922507964546621512713438470702986642486608412251521039 * 
--        97927786390663519429528993360368267006249228136794892056090651513080073109454331808866772457049032741774590681339704155886317906072752116837364369820881 * 
--        6311333012067573859934619875281580722169341118251824810685189958869028563705791257098179568281267604475713194506701767181158922314632507024334758203314465 , 
--        6703903964971298549787012499102923063739682910296196688861780721860882015036773488400937149083451713845015929093243025426876941405973284973216824503042159 ) = 
--        = 5770539552593938046267215339235143056108840937616962443047031076129629580294766891795665005337423591502330655021878623252853392851503861478061794255888635
--    where 6311333012067573859934619875281580722169341118251824810685189958869028563705791257098179568281267604475713194506701767181158922314632507024334758203314465 is the inverse modulus
--------------------------------------------------	  

      --    A = 3351951982485649274893506249551461531869841455148098344430890360930441007518386744200468574541725856922507964546621512713438470702986642486608412251521039 in decimal
      A <=  "01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111";
      --    B = 97927786390663519429528993360368267006249228136794892056090651513080073109454331808866772457049032741774590681339704155886317906072752116837364369820881 in decimal
	  B <=  "00000001110111101010100100111010100000100100111111101001100100111011001111000010101011111001001001110011011010010100101000100010110011011101111000010011100100101000011010000110110010101101101100000111101000001111010101000110100001100011101110100011100111101100000001000110010110111001110111111110101000001110001000011001000001000000111100000001100110000100011100010011101110010100111110010111110001000110111010010010101101001111110000111001110000100111111111100011011101100000011110100100100000011000110011010001";
      --    M = 6703903964971298549787012499102923063739682910296196688861780721860882015036773488400937149083451713845015929093243025426876941405973284973216824503042159 in decimal
      M <=  "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111";
		wait for clk_period;
--    Result = 1075674849379283795 in decimal	
		start <= '1';
		
		--wait for 600*clk_period;
		wait until ready = '1' and clk = '0';
	  if product /= x"6e2dcf4e2226cb7a14afa007b0bafdf50d573776681c0cca8d7ff56515076baffd05eaa8ee73d63874a1df6d13e2bbc0aeb6dcd21d8ee10613df1e2e5e02e0fb" then
        report "RESULT MISMATCH! Test case 2 failed" severity ERROR;
		assert false severity failure;
	  else
		report "Test case 2 successful" severity note;	
	  end if; 
		
		assert false severity failure;
   end process;

END;
