--------------------------------------------------------------------------------
-- Company: 
--
-- File: cp_FullAdder.vhd
--
-- Description:
--	projet copyblaze
--	1 bit Full adder
--
-- File history:
-- v1.0: 14/10/11: Creation
--
-- Targeted device: ProAsic A3P250 VQFP100
-- Author: AbdAllah Meziti
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use	work.Usefull_Pkg.all;		-- Usefull Package

--------------------------------------------------------------------------------
-- Entity: cp_FullAdder
--
-- Description:
--	
--	REMARQUE:
--
--	
-- History:
-- 14/10/11 AM: Creation
-- ---------------------
-- xx/xx/xx AM: 
--				
--------------------------------------------------------------------------------
entity cp_FullAdder is
	port (
	--------------------------------------------------------------------------------
	-- Signaux Fonctionels
	--------------------------------------------------------------------------------
		Ci_i		: in std_ulogic;
		A_i			: in std_ulogic;
		B_i			: in std_ulogic;

		Co_o		: out std_ulogic;
		S_o			: out std_ulogic
	);
end cp_FullAdder;

--------------------------------------------------------------------------------
-- Architecture: RTL
-- of entity : cp_FullAdder
--------------------------------------------------------------------------------
architecture rtl of cp_FullAdder is

	--------------------------------------------------------------------------------
	-- D�finition des fonctions
	--------------------------------------------------------------------------------
	


	--------------------------------------------------------------------------------
	-- D�finition des constantes
	--------------------------------------------------------------------------------

	--------------------------------------------------------------------------------
	-- D�finition des signaux interne
	--------------------------------------------------------------------------------

	--------------------------------------------------------------------------------
	-- D�claration des composants
	--------------------------------------------------------------------------------

begin

	--------------------------------------------------------------------------------
	-- Full adder
	--------------------------------------------------------------------------------
	-- SUM
	S_o		<=	A_i xor B_i xor Ci_i;
	-- CARRY
	Co_o	<=	(A_i and B_i) or (B_i and Ci_i) or (A_i and Ci_i);

end rtl;

