module Raptor64mc_tb();
parameter IDLE = 8'd1;
parameter DOCMD = 8'd2;

reg clk;
reg rst;
reg nmi;
wire sys_cyc;
wire sys_stb;
wire sys_we;
wire [7:0] sys_sel;
wire [31:0] sys_adr;
wire [31:0] sys_dbo;
wire [31:0] sys_dbi;
wire sys_ack;
wire cmd_en;
wire [2:0] cmd_instr;
wire [5:0] cmd_bl;
wire [29:0] cmd_byte_addr;
reg cmd_full;
reg [5:0] tb_cmd_bl;
reg [2:0] tb_cmd_instr;
reg [29:0] tb_cmd_byte_addr;
wire rd_en;
reg rd_empty;
reg [31:0] rd_data;
reg [7:0] cnt;
wire wr_en;
wire [31:0] wr_data;
wire wr_empty = 1'b1;
wire wr_full;
reg [31:0] iromout;

assign sys_ack = sys_stb;

initial begin
	clk = 1;
	rst = 0;
	nmi = 0;
	#100 rst = 1;
	#100 rst = 0;
	#1300 nmi = 1;
	#100 nmi = 0;
end

always #10 clk = ~clk;	//  50 MHz

always @(sys_adr)
case(sys_adr | 64'hFFFF_FFFF_FFFF_0000)
64'h70:	iromout <= 32'h00000020;
64'h74:	iromout <= 32'h00000000;
64'h78:	iromout <= 32'h000DE000;
64'h7C:	iromout <= 32'h37800000;
64'h80:	iromout <= 32'h00000000;
64'h84:	iromout <= 32'h00000378;
64'h88:	iromout <= 32'h000DE000;
64'h8C:	iromout <= 32'h37800000;
64'hFFFFFFFFFFFFF000:	iromout <= 32'h02000AA8;
64'hFFFFFFFFFFFFF004:	iromout <= 32'h00062408;
64'hFFFFFFFFFFFFF008:	iromout <= 32'h210BE100;
64'hFFFFFFFFFFFFF00C:	iromout <= 32'h0A176543;
64'hFFFFFFFFFFFFF010:	iromout <= 32'h400008A9;
64'hFFFFFFFFFFFFF014:	iromout <= 32'h0026A408;
64'hFFFFFFFFFFFFF018:	iromout <= 32'hA9802100;
64'hFFFFFFFFFFFFF01C:	iromout <= 32'h0A1FEDCB;
64'hFFFFFFFFFFFFF020:	iromout <= 32'h40000929;
64'hFFFFFFFFFFFFF024:	iromout <= 32'h0028A408;
64'hFFFFFFFFFFFFF028:	iromout <= 32'h08802100;
64'hFFFFFFFFFFFFF02C:	iromout <= 32'h2F800000;
64'hFFFFFFFFFFFFF030:	iromout <= 32'h020013FD;
64'hFFFFFFFFFFFFF034:	iromout <= 32'h0010AC58;
64'hFFFFFFFFFFFFF038:	iromout <= 32'h01816010;
64'hFFFFFFFFFFFFF03C:	iromout <= 32'h01044500;
64'hFFFFFFFFFFFFF040:	iromout <= 32'hFFFFFFFF;
64'hFFFFFFFFFFFFF044:	iromout <= 32'h400003FF;
64'hFFFFFFFFFFFFF048:	iromout <= 32'h0321600F;
64'hFFFFFFFFFFFFF04C:	iromout <= 32'h05804000;
64'hFFFFFFFFFFFFF050:	iromout <= 32'h06000014;
64'hFFFFFFFFFFFFF054:	iromout <= 32'h00000058;
64'hFFFFFFFFFFFFF058:	iromout <= 32'h00262110;
64'hFFFFFFFFFFFFF05C:	iromout <= 32'h02842000;
64'hFFFFFFFFFFFFF060:	iromout <= 32'hC6000001;
64'hFFFFFFFFFFFFF064:	iromout <= 32'hFFFEA430;
64'hFFFFFFFFFFFFF068:	iromout <= 32'hC24BE307;
64'hFFFFFFFFFFFFF06C:	iromout <= 32'h0C7FFFFF;
64'hFFFFFFFFFFFFF070:	iromout <= 32'h00000000;
64'hFFFFFFFFFFFFF074:	iromout <= 32'h00000378;
64'hFFFFFFFFFFFFF078:	iromout <= 32'h000DE000;
64'hFFFFFFFFFFFFF07C:	iromout <= 32'h37800000;
64'hFFFFFFFFFFFFF090:	iromout <= 32'hFFFFFFFF;
64'hFFFFFFFFFFFFF094:	iromout <= 32'h700003FF;
64'hFFFFFFFFFFFFF098:	iromout <= 32'h0001600F;
64'hFFFFFFFFFFFFF09C:	iromout <= 32'h10044000;
64'hFFFFFFFFFFFFF0A0:	iromout <= 32'h81FFFFC1;
64'hFFFFFFFFFFFFF0A4:	iromout <= 32'h000006F8;
64'hFFFFFFFFFFFFF0A8:	iromout <= 32'h00040100;
64'hFFFFFFFFFFFFF0AC:	iromout <= 32'h0D83E000;
64'hFFFFFFFFFFFFF0B0:	iromout <= 32'h00800009;
64'hFFFFFFFFFFFFF0B4:	iromout <= 32'hAAAB5410;
64'hFFFFFFFFFFFFF0B8:	iromout <= 32'h555F5554;
64'hFFFFFFFFFFFFF0BC:	iromout <= 32'h05802AA5;
64'hFFFFFFFFFFFFF0C0:	iromout <= 32'h02000000;
64'hFFFFFFFFFFFFF0C4:	iromout <= 32'h0000019A;
64'hFFFFFFFFFFFFF0C8:	iromout <= 32'h00646810;
64'hFFFFFFFFFFFFF0CC:	iromout <= 32'h01044300;
64'hFFFFFFFFFFFFF0D0:	iromout <= 32'hC00000A9;
64'hFFFFFFFFFFFFF0D4:	iromout <= 32'h000022F8;
64'hFFFFFFFFFFFFF0D8:	iromout <= 32'h0000A840;
64'hFFFFFFFFFFFFF0DC:	iromout <= 32'h04206000;
64'hFFFFFFFFFFFFF0E0:	iromout <= 32'hC1FFFF00;
64'hFFFFFFFFFFFFF0E4:	iromout <= 32'h800026F8;
64'hFFFFFFFFFFFFF0E8:	iromout <= 32'h00904802;
64'hFFFFFFFFFFFFF0EC:	iromout <= 32'h01000800;
64'hFFFFFFFFFFFFF0F0:	iromout <= 32'h04000000;
64'hFFFFFFFFFFFFF0F4:	iromout <= 32'hA955551A;
64'hFFFFFFFFFFFFF0F8:	iromout <= 32'h1091021A;
64'hFFFFFFFFFFFFF0FC:	iromout <= 32'h2F8C0000;
64'hFFFFFFFFFFFFF100:	iromout <= 32'h10000008;
64'hFFFFFFFFFFFFF104:	iromout <= 32'h00000022;
64'hFFFFFFFFFFFFF108:	iromout <= 32'hF801081C;
64'hFFFFFFFFFFFFF10C:	iromout <= 32'h2F8C1FFF;
64'hFFFFFFFFFFFFF110:	iromout <= 32'h14000329;
64'hFFFFFFFFFFFFF114:	iromout <= 32'h000026FA;
64'hFFFFFFFFFFFFF118:	iromout <= 32'h52A04002;
64'hFFFFFFFFFFFFF11C:	iromout <= 32'h3AAAAD55;
64'hFFFFFFFFFFFFF120:	iromout <= 32'h0355AAAA;
64'hFFFFFFFFFFFFF124:	iromout <= 32'h00000058;
64'hFFFFFFFFFFFFF128:	iromout <= 32'h00066808;
64'hFFFFFFFFFFFFF12C:	iromout <= 32'h11A04000;
64'hFFFFFFFFFFFFF130:	iromout <= 32'h44300006;
64'hFFFFFFFFFFFFF134:	iromout <= 32'h00032410;
64'hFFFFFFFFFFFFF138:	iromout <= 32'h008BE300;
64'hFFFFFFFFFFFFF13C:	iromout <= 32'h02210000;
64'hFFFFFFFFFFFFF140:	iromout <= 32'h07000000;
64'hFFFFFFFFFFFFF144:	iromout <= 32'hFFFC8042;
64'hFFFFFFFFFFFFF148:	iromout <= 32'h009BE307;
64'hFFFFFFFFFFFFF14C:	iromout <= 32'h01200B00;
64'hFFFFFFFFFFFFF150:	iromout <= 32'h00800009;
64'hFFFFFFFFFFFFF154:	iromout <= 32'h00000010;
64'hFFFFFFFFFFFFF158:	iromout <= 32'hAAA46810;
64'hFFFFFFFFFFFFF15C:	iromout <= 32'h0408755A;
64'hFFFFFFFFFFFFF160:	iromout <= 32'hC00000A9;
64'hFFFFFFFFFFFFF164:	iromout <= 32'h000022F8;
64'hFFFFFFFFFFFFF168:	iromout <= 32'h00008840;
64'hFFFFFFFFFFFFF16C:	iromout <= 32'h04207000;
64'hFFFFFFFFFFFFF170:	iromout <= 32'hC1FFFF20;
64'hFFFFFFFFFFFFF174:	iromout <= 32'h000222F8;
64'hFFFFFFFFFFFFF178:	iromout <= 32'h014BE858;
64'hFFFFFFFFFFFFF17C:	iromout <= 32'h01216800;
64'hFFFFFFFFFFFFF180:	iromout <= 32'h14000048;
64'hFFFFFFFFFFFFF184:	iromout <= 32'h000052FA;
64'hFFFFFFFFFFFFF188:	iromout <= 32'h40004852;
64'hFFFFFFFFFFFFF18C:	iromout <= 32'h19810000;
64'hFFFFFFFFFFFFF190:	iromout <= 32'h3E000000;
64'hFFFFFFFFFFFFF194:	iromout <= 32'h000080D8;
64'hFFFFFFFFFFFFF198:	iromout <= 32'h03400000;
64'hFFFFFFFFFFFFF19C:	iromout <= 32'h00802000;
64'hFFFFFFFFFFFFF1A0:	iromout <= 32'h41FFFFC9;
64'hFFFFFFFFFFFFF1A4:	iromout <= 32'hFC0002F8;
64'hFFFFFFFFFFFFF1A8:	iromout <= 32'h0086600F;
64'hFFFFFFFFFFFFF1AC:	iromout <= 32'h19805FF0;
64'hFFFFFFFFFFFFF1B0:	iromout <= 32'h02000228;
64'hFFFFFFFFFFFFF1B4:	iromout <= 32'h0010A008;
64'hFFFFFFFFFFFFF1B8:	iromout <= 32'hFA902010;
64'hFFFFFFFFFFFFF1BC:	iromout <= 32'hFFFFFFFF;
64'hFFFFFFFFFFFFF1C0:	iromout <= 32'h84680001;
64'hFFFFFFFFFFFFF1C4:	iromout <= 32'h40000C18;
64'hFFFFFFFFFFFFF1C8:	iromout <= 32'h00004110;
64'hFFFFFFFFFFFFF1CC:	iromout <= 32'h11844000;
64'hFFFFFFFFFFFFF1D0:	iromout <= 32'hFFFFFFA9;
64'hFFFFFFFFFFFFF1D4:	iromout <= 32'h0000CFFF;
64'hFFFFFFFFFFFFF1D8:	iromout <= 32'h03502000;
64'hFFFFFFFFFFFFF1DC:	iromout <= 32'h00800000;
64'hFFFFFFFFFFFFF1E0:	iromout <= 32'h03FF0000;
64'hFFFFFFFFFFFFF1E4:	iromout <= 32'hFC002118;
64'hFFFFFFFFFFFFF1E8:	iromout <= 32'h02046017;
64'hFFFFFFFFFFFFF1EC:	iromout <= 32'h00000000;
64'hFFFFFFFFFFFFFFB0:	iromout <= 32'hFFFFFC66;
64'hFFFFFFFFFFFFFFB4:	iromout <= 32'h000000CF;
64'hFFFFFFFFFFFFFFB8:	iromout <= 32'h000DE000;
64'hFFFFFFFFFFFFFFBC:	iromout <= 32'h37800000;
64'hFFFFFFFFFFFFFFC0:	iromout <= 32'hFFFFFC66;
64'hFFFFFFFFFFFFFFC4:	iromout <= 32'h000000CF;
64'hFFFFFFFFFFFFFFC8:	iromout <= 32'h000DE000;
64'hFFFFFFFFFFFFFFCC:	iromout <= 32'h37800000;
64'hFFFFFFFFFFFFFFD0:	iromout <= 32'h00000000;
64'hFFFFFFFFFFFFFFD4:	iromout <= 32'h00000378;
64'hFFFFFFFFFFFFFFD8:	iromout <= 32'h000DE000;
64'hFFFFFFFFFFFFFFDC:	iromout <= 32'h37800000;
64'hFFFFFFFFFFFFFFE0:	iromout <= 32'hFFFFFC65;
64'hFFFFFFFFFFFFFFE4:	iromout <= 32'h000000CF;
64'hFFFFFFFFFFFFFFE8:	iromout <= 32'h000DE000;
64'hFFFFFFFFFFFFFFEC:	iromout <= 32'h37800000;
64'hFFFFFFFFFFFFFFF0:	iromout <= 32'hFFFFFC00;
64'hFFFFFFFFFFFFFFF4:	iromout <= 32'h000000CF;
64'hFFFFFFFFFFFFFFF8:	iromout <= 32'h00000000;
64'hFFFFFFFFFFFFFFFC:	iromout <= 32'h00000000;
endcase
assign sys_dbi = iromout;

reg [7:0] state;
always @(posedge clk)
if (rst) begin
	state <= IDLE;
	cmd_full <= 1'b0;
	rd_empty <= 1'b1;
end
else begin
case(state)
IDLE:
	if (cmd_en) begin
		tb_cmd_instr <= cmd_instr;
		tb_cmd_bl <= cmd_bl;
		tb_cmd_byte_addr <= cmd_byte_addr;
		cmd_full <= 1'b1;
		rd_empty <= 1'b1;
		cnt <= 8'd0;
		state <= DOCMD;
	end
DOCMD:
	case(tb_cmd_instr)
	3'b000:	
		begin
			cmd_full <= 1'b0;
			state <= IDLE;
		end
	2'b001:
		begin
			cmd_full <= 1'b0;
			state <= IDLE;
		end
	endcase
default:	state <= IDLE;
endcase
	if (rd_en) begin
		if (cnt>=3) begin
			rd_empty <= 1'b0;
		case(tb_cmd_byte_addr | 64'hFFFF_FFFF_FFFF_0000)
64'hFFFFFFFFFFFFF000:	rd_data <= 32'h020013FD;
64'hFFFFFFFFFFFFF004:	rd_data <= 32'h00006050;
64'hFFFFFFFFFFFFF008:	rd_data <= 32'h01802120;
64'hFFFFFFFFFFFFF00C:	rd_data <= 32'h00848000;
64'hFFFFFFFFFFFFF010:	rd_data <= 32'h0400042B;
64'hFFFFFFFFFFFFF014:	rd_data <= 32'h40006050;
64'hFFFFFFFFFFFFF018:	rd_data <= 32'hFFF04111;
64'hFFFFFFFFFFFFF01C:	rd_data <= 32'h3FFFFFFF;
64'hFFFFFFFFFFFFF020:	rd_data <= 32'h03D00000;
64'hFFFFFFFFFFFFF024:	rd_data <= 32'h0000C850;
64'hFFFFFFFFFFFFF028:	rd_data <= 32'h64C14010;
64'hFFFFFFFFFFFFF02C:	rd_data <= 32'h05006000;
64'hFFFFFFFFFFFFF030:	rd_data <= 32'h44000000;
64'hFFFFFFFFFFFFF034:	rd_data <= 32'h00000988;
64'hFFFFFFFFFFFFF038:	rd_data <= 32'h0010A108;
64'hFFFFFFFFFFFFF03C:	rd_data <= 32'h030C6000;
64'hFFFFFFFFFFFFF040:	rd_data <= 32'hC1FFFF81;
64'hFFFFFFFFFFFFF044:	rd_data <= 32'hFFF062F8;
64'hFFFFFFFFFFFFF048:	rd_data <= 32'h00031FFF;
64'hFFFFFFFFFFFFF04C:	rd_data <= 32'h37800000;
64'hFFFFFFFFFFFFF050:	rd_data <= 32'h00000000;
64'hFFFFFFFFFFFFF054:	rd_data <= 32'h00000378;
64'hFFFFFFFFFFFFF058:	rd_data <= 32'h000DE000;
64'hFFFFFFFFFFFFF05C:	rd_data <= 32'h37800000;
64'hFFFFFFFFFFFFF060:	rd_data <= 32'hFFFFFFFF;
64'hFFFFFFFFFFFFF064:	rd_data <= 32'h700003FF;
64'hFFFFFFFFFFFFF068:	rd_data <= 32'h0001400F;
64'hFFFFFFFFFFFFF06C:	rd_data <= 32'h10044000;
64'hFFFFFFFFFFFFF070:	rd_data <= 32'h81FFFFC5;
64'hFFFFFFFFFFFFF074:	rd_data <= 32'h000006F8;
64'hFFFFFFFFFFFFF078:	rd_data <= 32'h00040100;
64'hFFFFFFFFFFFFF07C:	rd_data <= 32'h0D83E000;
64'hFFFFFFFFFFFFF080:	rd_data <= 32'h00800009;
64'hFFFFFFFFFFFFF084:	rd_data <= 32'hAAAB5410;
64'hFFFFFFFFFFFFF088:	rd_data <= 32'h555F5554;
64'hFFFFFFFFFFFFF08C:	rd_data <= 32'h05002AA5;
64'hFFFFFFFFFFFFF090:	rd_data <= 32'h02000000;
64'hFFFFFFFFFFFFF094:	rd_data <= 32'h0000019A;
64'hFFFFFFFFFFFFF098:	rd_data <= 32'h00646810;
64'hFFFFFFFFFFFFF09C:	rd_data <= 32'h01044300;
64'hFFFFFFFFFFFFF0A0:	rd_data <= 32'hC00000A1;
64'hFFFFFFFFFFFFF0A4:	rd_data <= 32'h000022F8;
64'hFFFFFFFFFFFFF0A8:	rd_data <= 32'h0000A840;
64'hFFFFFFFFFFFFF0AC:	rd_data <= 32'h03A06000;
64'hFFFFFFFFFFFFF0B0:	rd_data <= 32'hC1FFFF02;
64'hFFFFFFFFFFFFF0B4:	rd_data <= 32'h800026F8;
64'hFFFFFFFFFFFFF0B8:	rd_data <= 32'h00904802;
64'hFFFFFFFFFFFFF0BC:	rd_data <= 32'h01000800;
64'hFFFFFFFFFFFFF0C0:	rd_data <= 32'h04000000;
64'hFFFFFFFFFFFFF0C4:	rd_data <= 32'hA955551A;
64'hFFFFFFFFFFFFF0C8:	rd_data <= 32'h1010E21A;
64'hFFFFFFFFFFFFF0CC:	rd_data <= 32'h2F8C0000;
64'hFFFFFFFFFFFFF0D0:	rd_data <= 32'h10000008;
64'hFFFFFFFFFFFFF0D4:	rd_data <= 32'h00000022;
64'hFFFFFFFFFFFFF0D8:	rd_data <= 32'hF820E81C;
64'hFFFFFFFFFFFFF0DC:	rd_data <= 32'h2F8C1FFF;
64'hFFFFFFFFFFFFF0E0:	rd_data <= 32'h14000321;
64'hFFFFFFFFFFFFF0E4:	rd_data <= 32'h000026FA;
64'hFFFFFFFFFFFFF0E8:	rd_data <= 32'h52A04002;
64'hFFFFFFFFFFFFF0EC:	rd_data <= 32'h3AAAAD55;
64'hFFFFFFFFFFFFF0F0:	rd_data <= 32'h0355AAAA;
64'hFFFFFFFFFFFFF0F4:	rd_data <= 32'h00000050;
64'hFFFFFFFFFFFFF0F8:	rd_data <= 32'h00066808;
64'hFFFFFFFFFFFFF0FC:	rd_data <= 32'h11A04000;
64'hFFFFFFFFFFFFF100:	rd_data <= 32'h44300006;
64'hFFFFFFFFFFFFF104:	rd_data <= 32'h00030410;
64'hFFFFFFFFFFFFF108:	rd_data <= 32'h008BE300;
64'hFFFFFFFFFFFFF10C:	rd_data <= 32'h02210000;
64'hFFFFFFFFFFFFF110:	rd_data <= 32'h07000000;
64'hFFFFFFFFFFFFF114:	rd_data <= 32'hFFFC883A;
64'hFFFFFFFFFFFFF118:	rd_data <= 32'h009BE307;
64'hFFFFFFFFFFFFF11C:	rd_data <= 32'h01200B00;
64'hFFFFFFFFFFFFF120:	rd_data <= 32'h00800009;
64'hFFFFFFFFFFFFF124:	rd_data <= 32'h00000010;
64'hFFFFFFFFFFFFF128:	rd_data <= 32'hAAA46810;
64'hFFFFFFFFFFFFF12C:	rd_data <= 32'h0388755A;
64'hFFFFFFFFFFFFF130:	rd_data <= 32'hC00000A1;
64'hFFFFFFFFFFFFF134:	rd_data <= 32'h000022F8;
64'hFFFFFFFFFFFFF138:	rd_data <= 32'h00008840;
64'hFFFFFFFFFFFFF13C:	rd_data <= 32'h03A07000;
64'hFFFFFFFFFFFFF140:	rd_data <= 32'hC1FFFF22;
64'hFFFFFFFFFFFFF144:	rd_data <= 32'h000202F8;
64'hFFFFFFFFFFFFF148:	rd_data <= 32'h014BE858;
64'hFFFFFFFFFFFFF14C:	rd_data <= 32'h01216800;
64'hFFFFFFFFFFFFF150:	rd_data <= 32'h14000040;
64'hFFFFFFFFFFFFF154:	rd_data <= 32'h000052FA;
64'hFFFFFFFFFFFFF158:	rd_data <= 32'h40004852;
64'hFFFFFFFFFFFFF15C:	rd_data <= 32'h19810000;
64'hFFFFFFFFFFFFF160:	rd_data <= 32'h3E000000;
64'hFFFFFFFFFFFFF164:	rd_data <= 32'h0000C8D8;
64'hFFFFFFFFFFFFF168:	rd_data <= 32'h02102008;
64'hFFFFFFFFFFFFF16C:	rd_data <= 32'h2F840000;
64'hFFFFFFFFFFFFF170:	rd_data <= 32'h03FF0000;
64'hFFFFFFFFFFFFF174:	rd_data <= 32'hFC002198;
64'hFFFFFFFFFFFFF178:	rd_data <= 32'h22866017;
64'hFFFFFFFFFFFFF17C:	rd_data <= 32'h00802000;
64'hFFFFFFFFFFFFF180:	rd_data <= 32'h04000428;
64'hFFFFFFFFFFFFF184:	rd_data <= 32'h0016A408;
64'hFFFFFFFFFFFFF188:	rd_data <= 32'h00102200;
64'hFFFFFFFFFFFFF18C:	rd_data <= 32'h01884680;
64'hFFFFFFFFFFFFF190:	rd_data <= 32'h44100003;
64'hFFFFFFFFFFFFF194:	rd_data <= 32'h00000010;
64'hFFFFFFFFFFFFF198:	rd_data <= 32'h52946110;
64'hFFFFFFFFFFFFF19C:	rd_data <= 32'h00880000;
64'hFFFFFFFFFFFFF1A0:	rd_data <= 32'h00000034;
64'hFFFFFFFFFFFFF1A4:	rd_data <= 32'h0000CC08;
64'hFFFFFFFFFFFFF1A8:	rd_data <= 32'h00002000;
64'hFFFFFFFFFFFFF1AC:	rd_data <= 32'h11803FF0;
64'hFFFFFFFFFFFFF1B0:	rd_data <= 32'h05FF0008;
64'hFFFFFFFFFFFFF1B4:	rd_data <= 32'h00008118;
64'hFFFFFFFFFFFFF1B8:	rd_data <= 32'h00000000;
64'hFFFFFFFFFFFFF1BC:	rd_data <= 32'h37800000;
64'hFFFFFFFFFFFFFFB0:	rd_data <= 32'hFFFFFC59;
64'hFFFFFFFFFFFFFFB4:	rd_data <= 32'h000000CF;
64'hFFFFFFFFFFFFFFB8:	rd_data <= 32'h000DE000;
64'hFFFFFFFFFFFFFFBC:	rd_data <= 32'h37800000;
64'hFFFFFFFFFFFFFFC0:	rd_data <= 32'h00000000;
64'hFFFFFFFFFFFFFFC4:	rd_data <= 32'h00000378;
64'hFFFFFFFFFFFFFFC8:	rd_data <= 32'h000DE000;
64'hFFFFFFFFFFFFFFCC:	rd_data <= 32'h37800000;
64'hFFFFFFFFFFFFFFD0:	rd_data <= 32'h00000000;
64'hFFFFFFFFFFFFFFD4:	rd_data <= 32'h00000378;
64'hFFFFFFFFFFFFFFD8:	rd_data <= 32'h000DE000;
64'hFFFFFFFFFFFFFFDC:	rd_data <= 32'h37800000;
64'hFFFFFFFFFFFFFFE0:	rd_data <= 32'h00000000;
64'hFFFFFFFFFFFFFFE4:	rd_data <= 32'h00000378;
64'hFFFFFFFFFFFFFFE8:	rd_data <= 32'h000DE000;
64'hFFFFFFFFFFFFFFEC:	rd_data <= 32'h37800000;
64'hFFFFFFFFFFFFFFF0:	rd_data <= 32'hFFFFFC00;
64'hFFFFFFFFFFFFFFF4:	rd_data <= 32'h000000CF;
64'hFFFFFFFFFFFFFFF8:	rd_data <= 32'h00000000;
64'hFFFFFFFFFFFFFFFC:	rd_data <= 32'h00000000;

//		30'h0:	rd_data <= 32'h00000000;
//		30'h4:	rd_data <= 32'h00002378;
//		30'h8:	rd_data <= 32'h00030000;
//		30'hC:	rd_data <= 32'h37800000;
//		30'h10:	rd_data <= 32'h00000000;
//		30'h14:	rd_data <= 32'h00000378;
//		30'h18:	rd_data <= 32'h000DE000;
//		30'h1C:	rd_data <= 32'h37800000;
//		30'h20:	rd_data <= 32'hFFFFFFFF;
//		30'h24:	rd_data <= 32'h700003FF;
//		30'h28:	rd_data <= 32'h0001200F;
//		30'h2C:	rd_data <= 32'h0D83E000;
		endcase
		tb_cmd_byte_addr <= tb_cmd_byte_addr + 30'd4;
		tb_cmd_bl <= tb_cmd_bl - 6'd1;
		if (tb_cmd_bl==6'h0) rd_empty <= 1'b1;
		end
		else
			cnt <= cnt + 1;
	end
end

Raptor64mc u1
(
	.rst_i(rst),
	.clk_i(clk),
	.nmi_i(nmi),
	.irq_i(1'b0),
	.bte_o(),
	.cti_o(),
	.cyc_o(sys_cyc),
	.stb_o(sys_stb),
	.ack_i(sys_ack),
	.we_o(sys_we),
	.sel_o(sys_sel),
	.adr_o(sys_adr),
	.dat_i(sys_dbi),
	.dat_o(sys_dbo),

	.cmd_en(cmd_en),
	.cmd_instr(cmd_instr),
	.cmd_bl(cmd_bl),
	.cmd_byte_addr(cmd_byte_addr),
	.cmd_full(cmd_full),
	
	.rd_en(rd_en),
	.rd_data(rd_data),
	.rd_empty(rd_empty),

	.wr_en(wr_en),
	.wr_data(wr_data),
	.wr_full(1'b0),
	.wr_empty(1'b1),

	.sys_adv(1'b0),
	.sys_adr(59'd0)
);
endmodule
