//  #: Main
//  #: IP_PACKET
//  #: LAB_DAT
//  #: INI_DAT
//  #: BEG_DAT
//  #: END_DAT
//  #: LAB_ACK
//  #: LAB_CON
//  #: LAB_DRQ
//  #: DRQ_LOOP
//  #: END_DRQ
//  #: LAB_SENDACK
// labels:  {'DRQ_LOOP': 263, 'END_DRQ': 267, 'Main': 5, 'LAB_ACK': 161, 'LAB_SENDACK': 270, 'BEG_DAT': 153, 'LAB_DRQ': 190, 'LAB_CON': 168, 'INI_DAT': 149, 'LAB_DAT': 140, 'END_DAT': 157, 'IP_PACKET': 100}

module microcodesrc
(
	input		wire	[8:0]		addr,
	output	reg	[66:0]	code
);

always @(addr)
begin
	case (addr)

		// code: {	         <jmp,rst>
		//				         |      <in_rdy,out_rdy,aeof,asof>
		//				         |      |        <predmode>
		//				         |      |        |     <pred: fcs,eof,sof,equ,dst,src>
		//				         |      |        |     |          <High Byte Reg En>
		//				         |      |        |     |          |     <Output Byte Select>
		//				         |      |        |     |          |     |     <Outport_reg_en, Inport_eg_en>
		//				         |      |        |     |          |     |     |      <Data Mux Select>
		//				         |      |        |     |          |     |     |      |     <Op 0 Select>
		//				         |      |        |     |          |     |     |      |     |     <Op 1 Select>
		//				         |      |        |     |          |     |     |      |     |     |     <Register Address>
		//				         |      |        |     |          |     |     |      |     |     |     |       <Register Write Enables>
		//				         |      |        |     |          |     |     |      |     |     |     |       |     <FCS Add, FCS Clear>
		//				         |      |        |     |          |     |     |      |     |     |     |       |     |      <sr1ie,sr2ie,sr1oe,sr2oe>
		//				         |      |        |     |          |     |     |      |     |     |     |       |     |      |        <Flag Register>
		//				         |      |        |     |          |     |     |      |     |     |     |       |     |      |        |     <Compare Mode>
		//				         |      |        |     |          |     |     |      |     |     |     |       |     |      |        |     |     <ALU Op>
		//				         |      |        |     |          |     |     |      |     |     |     |       |     |      |        |     |     |     <Byte Constant>
		//				         |      |        |     |          |     |     |      |     |     |     |       |     |      |        |     |     |     |       <Word Constant> }
		000:			code <= {2'b10, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd1, 4'd10, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd1, 9'd005, 16'd00001}; // JMP(5, Cond=<IF: pred=[<<Constant: value=1>==<Register: address=10, high=True, low=True, high_byte_s=False>, Bytewide: False>]>, Flags=None)
		001:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd06, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // MOV(<Constant: value=0>,<Register: address=6, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		002:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd07, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // MOV(<Constant: value=0>,<Register: address=7, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		003:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd08, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // MOV(<Constant: value=0>,<Register: address=8, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		004:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd10, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // MOV(<Constant: value=1>,<Register: address=10, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		005:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b01, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // MOV(<Constant: value=0>,<Input Port Register>, Cond=None, Flags=None)
		006:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b10, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // MOV(<Constant: value=0>,<Output Port Register>, Cond=None, Flags=None)
		007:			code <= {2'b00, 4'b1000, 2'd1, 6'b001001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=<UNTIL: pred=[<SOF>, SRC]>, Flags=None)
		008:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		009:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		010:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		011:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		012:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		013:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		014:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		015:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		016:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		017:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		018:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		019:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		020:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Register: address=0, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		021:			code <= {2'b10, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd1, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd1, 9'd100, 16'd02048}; // JMP(100, Cond=<IF: pred=[<<Constant: value=2048>==<Register: address=0, high=True, low=True, high_byte_s=False>, Bytewide: False>]>, Flags=None)
		022:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd1, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd3, 2'd1, 9'd000, 16'd02054}; // RST(Cond=<IF: pred=[<<Constant: value=2054>!=<Register: address=0, high=True, low=True, high_byte_s=False>, Bytewide: False>]>, Flags=None)
		023:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		024:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		025:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		026:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Register: address=0, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		027:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd1, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd3, 2'd1, 9'd000, 16'd02048}; // RST(Cond=<IF: pred=[<<Constant: value=2048>!=<Register: address=0, high=True, low=True, high_byte_s=False>, Bytewide: False>]>, Flags=None)
		028:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		029:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		030:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		031:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Register: address=0, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		032:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd1, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd3, 2'd1, 9'd000, 16'd00001}; // RST(Cond=<IF: pred=[<<Constant: value=1>!=<Register: address=0, high=True, low=True, high_byte_s=False>, Bytewide: False>]>, Flags=None)
		033:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		034:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		035:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		036:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		037:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		038:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		039:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		040:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		041:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		042:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		043:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		044:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		045:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		046:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		047:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		048:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		049:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd7, 2'd1, 9'd000, 16'd00010}; // RST(Cond=<IF: pred=[<<Port>!=<Constant: value=10>, Bytewide: True>]>, Flags=None)
		050:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		051:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd7, 2'd1, 9'd000, 16'd00000}; // RST(Cond=<IF: pred=[<<Port>!=<Constant: value=0>, Bytewide: True>]>, Flags=None)
		052:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		053:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd7, 2'd1, 9'd000, 16'd00001}; // RST(Cond=<IF: pred=[<<Port>!=<Constant: value=1>, Bytewide: True>]>, Flags=None)
		054:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		055:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd7, 2'd1, 9'd000, 16'd00042}; // RST(Cond=<IF: pred=[<<Port>!=<Constant: value=42>, Bytewide: True>]>, Flags=None)
		056:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		057:			code <= {2'b00, 4'b0110, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=[<ASOF>])
		058:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		059:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		060:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		061:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		062:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		063:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // OUT(<Constant: value=1>, Cond=None, Flags=None)
		064:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00035}; // OUT(<Constant: value=35>, Cond=None, Flags=None)
		065:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00069}; // OUT(<Constant: value=69>, Cond=None, Flags=None)
		066:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00103}; // OUT(<Constant: value=103>, Cond=None, Flags=None)
		067:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00137}; // OUT(<Constant: value=137>, Cond=None, Flags=None)
		068:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00171}; // OUT(<Constant: value=171>, Cond=None, Flags=None)
		069:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00008}; // OUT(<Constant: value=8>, Cond=None, Flags=None)
		070:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00006}; // OUT(<Constant: value=6>, Cond=None, Flags=None)
		071:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		072:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // OUT(<Constant: value=1>, Cond=None, Flags=None)
		073:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00008}; // OUT(<Constant: value=8>, Cond=None, Flags=None)
		074:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		075:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00006}; // OUT(<Constant: value=6>, Cond=None, Flags=None)
		076:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00004}; // OUT(<Constant: value=4>, Cond=None, Flags=None)
		077:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		078:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00002}; // OUT(<Constant: value=2>, Cond=None, Flags=None)
		079:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // OUT(<Constant: value=1>, Cond=None, Flags=None)
		080:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00035}; // OUT(<Constant: value=35>, Cond=None, Flags=None)
		081:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00069}; // OUT(<Constant: value=69>, Cond=None, Flags=None)
		082:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00103}; // OUT(<Constant: value=103>, Cond=None, Flags=None)
		083:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00137}; // OUT(<Constant: value=137>, Cond=None, Flags=None)
		084:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00171}; // OUT(<Constant: value=171>, Cond=None, Flags=None)
		085:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00010}; // OUT(<Constant: value=10>, Cond=None, Flags=None)
		086:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		087:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // OUT(<Constant: value=1>, Cond=None, Flags=None)
		088:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00042}; // OUT(<Constant: value=42>, Cond=None, Flags=None)
		089:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		090:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		091:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		092:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		093:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		094:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		095:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		096:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		097:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		098:			code <= {2'b00, 4'b0101, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=[<AEOF>])
		099:			code <= {2'b01, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // RST(Cond=None, Flags=None)
		100:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		101:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		102:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		103:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		104:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		105:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		106:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		107:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		108:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		109:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd7, 2'd1, 9'd000, 16'd00017}; // RST(Cond=<IF: pred=[<<Port>!=<Constant: value=17>, Bytewide: True>]>, Flags=None)
		110:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		111:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		112:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		113:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		114:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		115:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		116:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		117:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd7, 2'd1, 9'd000, 16'd00010}; // RST(Cond=<IF: pred=[<<Port>!=<Constant: value=10>, Bytewide: True>]>, Flags=None)
		118:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		119:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd7, 2'd1, 9'd000, 16'd00000}; // RST(Cond=<IF: pred=[<<Port>!=<Constant: value=0>, Bytewide: True>]>, Flags=None)
		120:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		121:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd7, 2'd1, 9'd000, 16'd00001}; // RST(Cond=<IF: pred=[<<Port>!=<Constant: value=1>, Bytewide: True>]>, Flags=None)
		122:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		123:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd7, 2'd1, 9'd000, 16'd00042}; // RST(Cond=<IF: pred=[<<Port>!=<Constant: value=42>, Bytewide: True>]>, Flags=None)
		124:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		125:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		126:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b1000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		127:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		128:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd3, 2'd1, 9'd000, 16'd12289}; // RST(Cond=<IF: pred=[<<Port>!=<Constant: value=12289>, Bytewide: False>]>, Flags=None)
		129:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		130:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		131:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		132:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		133:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		134:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Register: address=0, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		135:			code <= {2'b10, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd1, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd4, 2'd1, 9'd140, 16'd00000}; // JMP(140, Cond=<IF: pred=[<<Constant: value=0>==<Register: address=0, high=True, low=True, high_byte_s=False>, Bytewide: True>]>, Flags=None)
		136:			code <= {2'b10, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd1, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd4, 2'd1, 9'd161, 16'd00001}; // JMP(161, Cond=<IF: pred=[<<Constant: value=1>==<Register: address=0, high=True, low=True, high_byte_s=False>, Bytewide: True>]>, Flags=None)
		137:			code <= {2'b10, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd1, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd4, 2'd1, 9'd168, 16'd00002}; // JMP(168, Cond=<IF: pred=[<<Constant: value=2>==<Register: address=0, high=True, low=True, high_byte_s=False>, Bytewide: True>]>, Flags=None)
		138:			code <= {2'b10, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd1, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd4, 2'd1, 9'd190, 16'd00004}; // JMP(190, Cond=<IF: pred=[<<Constant: value=4>==<Register: address=0, high=True, low=True, high_byte_s=False>, Bytewide: True>]>, Flags=None)
		139:			code <= {2'b01, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // RST(Cond=None, Flags=None)
		140:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd09, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Register: address=9, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		141:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		142:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd1, 4'd06, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd3, 2'd1, 9'd000, 16'd00000}; // RST(Cond=<IF: pred=[<<Port>!=<Register: address=6, high=True, low=True, high_byte_s=False>, Bytewide: False>]>, Flags=None)
		143:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		144:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		145:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Register: address=0, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		146:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b10, 3'd2, 2'd0, 1'd0, 4'd09, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // MOV(<Register: address=9, high=True, low=True, high_byte_s=False>,<Output Port Register>, Cond=None, Flags=None)
		147:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd5, 2'd3, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd1, 9'd000, 16'd00001}; // SUB(<Register: address=0, high=True, low=True, high_byte_s=False>, <Constant: value=1>, <Register: address=0, high=True, low=True, high_byte_s=False>, Cond=NoneFlags=None)
		148:			code <= {2'b10, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd3, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd1, 9'd157, 16'd00000}; // JMP(157, Cond=<IF: pred=[<<Register: address=0, high=True, low=True, high_byte_s=False>==<Constant: value=0>, Bytewide: False>]>, Flags=None)
		149:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0100, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=2>, Cond=None, Flags=None)
		150:			code <= {2'b00, 4'b0110, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0001, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=2>, Cond=None, Flags=[<ASOF>])
		151:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd5, 2'd3, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd1, 9'd000, 16'd00001}; // SUB(<Register: address=0, high=True, low=True, high_byte_s=False>, <Constant: value=1>, <Register: address=0, high=True, low=True, high_byte_s=False>, Cond=NoneFlags=None)
		152:			code <= {2'b10, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd3, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd1, 9'd157, 16'd00000}; // JMP(157, Cond=<IF: pred=[<<Register: address=0, high=True, low=True, high_byte_s=False>==<Constant: value=0>, Bytewide: False>]>, Flags=None)
		153:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0100, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=2>, Cond=None, Flags=None)
		154:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0001, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=2>, Cond=None, Flags=None)
		155:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd5, 2'd3, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd1, 9'd000, 16'd00001}; // SUB(<Register: address=0, high=True, low=True, high_byte_s=False>, <Constant: value=1>, <Register: address=0, high=True, low=True, high_byte_s=False>, Cond=NoneFlags=None)
		156:			code <= {2'b10, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd3, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd3, 2'd1, 9'd153, 16'd00000}; // JMP(153, Cond=<IF: pred=[<<Register: address=0, high=True, low=True, high_byte_s=False>!=<Constant: value=0>, Bytewide: False>]>, Flags=None)
		157:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0100, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=2>, Cond=None, Flags=None)
		158:			code <= {2'b00, 4'b0101, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0001, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=2>, Cond=None, Flags=[<AEOF>])
		159:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b10, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // MOV(<Constant: value=0>,<Output Port Register>, Cond=None, Flags=None)
		160:			code <= {2'b10, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd270, 16'd00000}; // JMP(270, Cond=None, Flags=None)
		161:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		162:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		163:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd08, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Register: address=8, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		164:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		165:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		166:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		167:			code <= {2'b01, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // RST(Cond=None, Flags=None)
		168:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		169:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		170:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		171:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		172:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		173:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd03, 2'd2, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=3, high=True, low=False, high_byte_s=False>
		174:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd03, 2'd1, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=3, high=False, low=True, high_byte_s=False>
		175:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd04, 2'd2, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=4, high=True, low=False, high_byte_s=False>
		176:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd04, 2'd1, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=4, high=False, low=True, high_byte_s=False>
		177:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd05, 2'd2, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=5, high=True, low=False, high_byte_s=False>
		178:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd05, 2'd1, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=5, high=False, low=True, high_byte_s=False>
		179:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd01, 2'd2, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=1, high=True, low=False, high_byte_s=False>
		180:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd01, 2'd1, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=1, high=False, low=True, high_byte_s=False>
		181:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd02, 2'd2, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=2, high=True, low=False, high_byte_s=False>
		182:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd02, 2'd1, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=2, high=False, low=True, high_byte_s=False>
		183:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd12, 2'd2, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=12, high=True, low=False, high_byte_s=False>
		184:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd12, 2'd1, 2'b00, 4'b1010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // Copy and Wrap SR:<Shif Register: sr_num=1> to R:<Register: address=12, high=False, low=True, high_byte_s=False>
		185:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd06, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // MOV(<Constant: value=0>,<Register: address=6, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		186:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd07, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // MOV(<Constant: value=0>,<Register: address=7, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		187:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd08, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // MOV(<Constant: value=0>,<Register: address=8, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		188:			code <= {2'b10, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd270, 16'd00000}; // JMP(270, Cond=None, Flags=None)
		189:			code <= {2'b01, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // RST(Cond=None, Flags=None)
		190:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd09, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Register: address=9, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		191:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		192:			code <= {2'b01, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd1, 1'd1, 4'd06, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd3, 2'd1, 9'd000, 16'd00000}; // RST(Cond=<IF: pred=[<<Port>!=<Register: address=6, high=True, low=True, high_byte_s=False>, Bytewide: False>]>, Flags=None)
		193:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		194:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b1, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<High Byte Register>, Cond=None, Flags=None)
		195:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Register: address=0, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		196:			code <= {2'b00, 4'b0110, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=[<ASOF>])
		197:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		198:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		199:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		200:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		201:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		202:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // OUT(<Constant: value=1>, Cond=None, Flags=None)
		203:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00035}; // OUT(<Constant: value=35>, Cond=None, Flags=None)
		204:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00069}; // OUT(<Constant: value=69>, Cond=None, Flags=None)
		205:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00103}; // OUT(<Constant: value=103>, Cond=None, Flags=None)
		206:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00137}; // OUT(<Constant: value=137>, Cond=None, Flags=None)
		207:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00171}; // OUT(<Constant: value=171>, Cond=None, Flags=None)
		208:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00008}; // OUT(<Constant: value=8>, Cond=None, Flags=None)
		209:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		210:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b01, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSC()
		211:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd17664}; // CSA(<Constant: value=17664>)
		212:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00069}; // OUT(<Constant: value=69>, Cond=None, Flags=None)
		213:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		214:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd5, 2'd0, 1'd1, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00034}; // ADD(<Constant: value=34>, <Register: address=0, high=True, low=True, high_byte_s=False>, <Register: address=0, high=True, low=True, high_byte_s=False>, Cond=NoneFlags=None)
		215:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSA(<Register: address=0, high=True, low=True, high_byte_s=False>)
		216:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd1, 2'b00, 3'd2, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Register: address=0, high=True, low=True, high_byte_s=True>, Cond=None, Flags=None)
		217:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Register: address=0, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		218:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd5, 2'd3, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd1, 9'd000, 16'd00034}; // SUB(<Register: address=0, high=True, low=True, high_byte_s=False>, <Constant: value=34>, <Register: address=0, high=True, low=True, high_byte_s=False>, Cond=NoneFlags=None)
		219:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		220:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		221:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		222:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		223:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd08209}; // CSA(<Constant: value=8209>)
		224:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00032}; // OUT(<Constant: value=32>, Cond=None, Flags=None)
		225:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00017}; // OUT(<Constant: value=17>, Cond=None, Flags=None)
		226:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd02560}; // CSA(<Constant: value=2560>)
		227:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00298}; // CSA(<Constant: value=298>)
		228:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd01, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSA(<Register: address=1, high=True, low=True, high_byte_s=False>)
		229:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd02, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSA(<Register: address=2, high=True, low=True, high_byte_s=False>)
		230:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd1, 2'b00, 3'd1, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Checksum: high_byte_s=True>, Cond=None, Flags=None)
		231:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd1, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Checksum: high_byte_s=False>, Cond=None, Flags=None)
		232:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00010}; // OUT(<Constant: value=10>, Cond=None, Flags=None)
		233:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		234:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // OUT(<Constant: value=1>, Cond=None, Flags=None)
		235:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00042}; // OUT(<Constant: value=42>, Cond=None, Flags=None)
		236:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		237:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		238:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		239:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		240:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b01, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSC()
		241:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd12289}; // CSA(<Constant: value=12289>)
		242:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd12, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSA(<Register: address=12, high=True, low=True, high_byte_s=False>)
		243:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00048}; // OUT(<Constant: value=48>, Cond=None, Flags=None)
		244:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // OUT(<Constant: value=1>, Cond=None, Flags=None)
		245:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		246:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		247:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd5, 2'd0, 1'd1, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00014}; // ADD(<Constant: value=14>, <Register: address=0, high=True, low=True, high_byte_s=False>, <Register: address=0, high=True, low=True, high_byte_s=False>, Cond=NoneFlags=None)
		248:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd1, 2'b00, 3'd2, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Register: address=0, high=True, low=True, high_byte_s=True>, Cond=None, Flags=None)
		249:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Register: address=0, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		250:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSA(<Register: address=0, high=True, low=True, high_byte_s=False>)
		251:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd5, 2'd3, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd1, 9'd000, 16'd00014}; // SUB(<Register: address=0, high=True, low=True, high_byte_s=False>, <Constant: value=14>, <Register: address=0, high=True, low=True, high_byte_s=False>, Cond=NoneFlags=None)
		252:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		253:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		254:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00005}; // OUT(<Constant: value=5>, Cond=None, Flags=None)
		255:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd09, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Register: address=9, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		256:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd1, 2'b00, 3'd2, 2'd0, 1'd0, 4'd06, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Register: address=6, high=True, low=True, high_byte_s=True>, Cond=None, Flags=None)
		257:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd06, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Register: address=6, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		258:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd5, 2'd0, 1'd1, 4'd06, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // ADD(<Constant: value=1>, <Register: address=6, high=True, low=True, high_byte_s=False>, <Register: address=6, high=True, low=True, high_byte_s=False>, Cond=NoneFlags=None)
		259:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd1, 2'b00, 3'd2, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Register: address=0, high=True, low=True, high_byte_s=True>, Cond=None, Flags=None)
		260:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Register: address=0, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		261:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b01, 3'd2, 2'd0, 1'd0, 4'd09, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // MOV(<Register: address=9, high=True, low=True, high_byte_s=False>,<Input Port Register>, Cond=None, Flags=None)
		262:			code <= {2'b10, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd3, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd1, 9'd267, 16'd00001}; // JMP(267, Cond=<IF: pred=[<<Register: address=0, high=True, low=True, high_byte_s=False>==<Constant: value=1>, Bytewide: False>]>, Flags=None)
		263:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0100, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=2>, Cond=None, Flags=None)
		264:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0001, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=2>, Cond=None, Flags=None)
		265:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd5, 2'd3, 1'd0, 4'd00, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd1, 9'd000, 16'd00001}; // SUB(<Register: address=0, high=True, low=True, high_byte_s=False>, <Constant: value=1>, <Register: address=0, high=True, low=True, high_byte_s=False>, Cond=NoneFlags=None)
		266:			code <= {2'b10, 4'b0000, 2'd2, 6'b000100, 1'b0, 1'd0, 2'b00, 3'd0, 2'd3, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd3, 2'd1, 9'd263, 16'd00001}; // JMP(263, Cond=<IF: pred=[<<Register: address=0, high=True, low=True, high_byte_s=False>!=<Constant: value=1>, Bytewide: False>]>, Flags=None)
		267:			code <= {2'b00, 4'b1000, 2'd0, 6'b000001, 1'b0, 1'd0, 2'b00, 3'd3, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0100, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // IN(<Shif Register: sr_num=2>, Cond=None, Flags=None)
		268:			code <= {2'b00, 4'b0101, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0001, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=2>, Cond=None, Flags=[<AEOF>])
		269:			code <= {2'b01, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // RST(Cond=None, Flags=None)
		270:			code <= {2'b00, 4'b0110, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=[<ASOF>])
		271:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		272:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		273:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		274:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		275:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		276:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // OUT(<Constant: value=1>, Cond=None, Flags=None)
		277:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00035}; // OUT(<Constant: value=35>, Cond=None, Flags=None)
		278:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00069}; // OUT(<Constant: value=69>, Cond=None, Flags=None)
		279:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00103}; // OUT(<Constant: value=103>, Cond=None, Flags=None)
		280:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00137}; // OUT(<Constant: value=137>, Cond=None, Flags=None)
		281:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00171}; // OUT(<Constant: value=171>, Cond=None, Flags=None)
		282:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00008}; // OUT(<Constant: value=8>, Cond=None, Flags=None)
		283:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		284:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b01, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSC()
		285:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd17664}; // CSA(<Constant: value=17664>)
		286:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00069}; // OUT(<Constant: value=69>, Cond=None, Flags=None)
		287:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		288:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00034}; // CSA(<Constant: value=34>)
		289:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		290:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00034}; // OUT(<Constant: value=34>, Cond=None, Flags=None)
		291:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		292:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		293:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		294:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		295:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd08209}; // CSA(<Constant: value=8209>)
		296:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00032}; // OUT(<Constant: value=32>, Cond=None, Flags=None)
		297:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00017}; // OUT(<Constant: value=17>, Cond=None, Flags=None)
		298:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd02560}; // CSA(<Constant: value=2560>)
		299:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00298}; // CSA(<Constant: value=298>)
		300:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd01, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSA(<Register: address=1, high=True, low=True, high_byte_s=False>)
		301:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd02, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSA(<Register: address=2, high=True, low=True, high_byte_s=False>)
		302:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd1, 2'b00, 3'd1, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Checksum: high_byte_s=True>, Cond=None, Flags=None)
		303:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd1, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Checksum: high_byte_s=False>, Cond=None, Flags=None)
		304:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00010}; // OUT(<Constant: value=10>, Cond=None, Flags=None)
		305:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		306:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // OUT(<Constant: value=1>, Cond=None, Flags=None)
		307:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00042}; // OUT(<Constant: value=42>, Cond=None, Flags=None)
		308:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		309:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		310:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		311:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		312:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00048}; // OUT(<Constant: value=48>, Cond=None, Flags=None)
		313:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // OUT(<Constant: value=1>, Cond=None, Flags=None)
		314:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b01, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSC()
		315:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd12289}; // CSA(<Constant: value=12289>)
		316:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd12, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // CSA(<Register: address=12, high=True, low=True, high_byte_s=False>)
		317:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		318:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd4, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0010, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Shif Register: sr_num=1>, Cond=None, Flags=None)
		319:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		320:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00014}; // OUT(<Constant: value=14>, Cond=None, Flags=None)
		321:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b10, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00006}; // CSA(<Constant: value=6>)
		322:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		323:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		324:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // OUT(<Constant: value=1>, Cond=None, Flags=None)
		325:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		326:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd1, 2'b00, 3'd2, 2'd0, 1'd0, 4'd06, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Register: address=6, high=True, low=True, high_byte_s=True>, Cond=None, Flags=None)
		327:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd2, 2'd0, 1'd0, 4'd06, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Register: address=6, high=True, low=True, high_byte_s=False>, Cond=None, Flags=None)
		328:			code <= {2'b00, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd5, 2'd0, 1'd1, 4'd06, 2'd3, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00001}; // ADD(<Constant: value=1>, <Register: address=6, high=True, low=True, high_byte_s=False>, <Register: address=6, high=True, low=True, high_byte_s=False>, Cond=NoneFlags=None)
		329:			code <= {2'b00, 4'b0100, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=None)
		330:			code <= {2'b00, 4'b0101, 2'd0, 6'b000010, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // OUT(<Constant: value=0>, Cond=None, Flags=[<AEOF>])
		331:			code <= {2'b01, 4'b0000, 2'd0, 6'b000000, 1'b0, 1'd0, 2'b00, 3'd0, 2'd0, 1'd0, 4'd00, 2'd0, 2'b00, 4'b0000, 1'b0, 3'd0, 2'd0, 9'd000, 16'd00000}; // RST(Cond=None, Flags=None)

	default: code <= 0;
	endcase
	
end
endmodule
